
--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/ccs_in_v1.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;

PACKAGE ccs_in_pkg_v1 IS

COMPONENT ccs_in_v1
  GENERIC (
    rscid    : INTEGER;
    width    : INTEGER
  );
  PORT (
    idat   : OUT std_logic_vector(width-1 DOWNTO 0);
    dat    : IN  std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

END ccs_in_pkg_v1;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY ccs_in_v1 IS
  GENERIC (
    rscid : INTEGER;
    width : INTEGER
  );
  PORT (
    idat  : OUT std_logic_vector(width-1 DOWNTO 0);
    dat   : IN  std_logic_vector(width-1 DOWNTO 0)
  );
END ccs_in_v1;

ARCHITECTURE beh OF ccs_in_v1 IS
BEGIN

  idat <= dat;

END beh;


--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/ccs_out_v1.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;

PACKAGE ccs_out_pkg_v1 IS

COMPONENT ccs_out_v1
  GENERIC (
    rscid    : INTEGER;
    width    : INTEGER
  );
  PORT (
    dat    : OUT std_logic_vector(width-1 DOWNTO 0);
    idat   : IN  std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

END ccs_out_pkg_v1;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY ccs_out_v1 IS
  GENERIC (
    rscid : INTEGER;
    width : INTEGER
  );
  PORT (
    dat   : OUT std_logic_vector(width-1 DOWNTO 0);
    idat  : IN  std_logic_vector(width-1 DOWNTO 0)
  );
END ccs_out_v1;

ARCHITECTURE beh OF ccs_out_v1 IS
BEGIN

  dat <= idat;

END beh;


--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
PACKAGE mgc_io_sync_pkg_v2 IS

COMPONENT mgc_io_sync_v2
  GENERIC (
    valid    : INTEGER RANGE 0 TO 1
  );
  PORT (
    ld       : IN    std_logic;
    lz       : OUT   std_logic
  );
END COMPONENT;

END mgc_io_sync_pkg_v2;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY mgc_io_sync_v2 IS
  GENERIC (
    valid    : INTEGER RANGE 0 TO 1
  );
  PORT (
    ld       : IN    std_logic;
    lz       : OUT   std_logic
  );
END mgc_io_sync_v2;

ARCHITECTURE beh OF mgc_io_sync_v2 IS
BEGIN

  lz <= ld;

END beh;


--------> ./rtl.vhdl 
-- ----------------------------------------------------------------------
--  HLS HDL:        VHDL Netlister
--  HLS Version:    10.5c/896140 Production Release
--  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
-- 
--  Generated by:   dss545@hansolo.poly.edu
--  Generated date: Wed Feb  3 19:34:26 2021
-- ----------------------------------------------------------------------

-- 
-- ------------------------------------------------------------------
--  Design Unit:    fir_core_core_fsm
--  FSM Module
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.ccs_out_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;


ENTITY fir_core_core_fsm IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    fsm_output : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    for_C_2_tr0 : IN STD_LOGIC
  );
END fir_core_core_fsm;

ARCHITECTURE v1 OF fir_core_core_fsm IS
  -- Default Constants

  -- FSM State Type Declaration for fir_core_core_fsm_1
  TYPE fir_core_core_fsm_1_ST IS (main_C_0, for_C_0, for_C_1, for_C_2, main_C_1);

  SIGNAL state_var : fir_core_core_fsm_1_ST;
  SIGNAL state_var_NS : fir_core_core_fsm_1_ST;

BEGIN
  fir_core_core_fsm_1 : PROCESS (for_C_2_tr0, state_var)
  BEGIN
    CASE state_var IS
      WHEN for_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010");
        state_var_NS <= for_C_1;
      WHEN for_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100");
        state_var_NS <= for_C_2;
      WHEN for_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000");
        IF ( for_C_2_tr0 = '1' ) THEN
          state_var_NS <= main_C_1;
        ELSE
          state_var_NS <= for_C_0;
        END IF;
      WHEN main_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000");
        state_var_NS <= main_C_0;
      -- main_C_0
      WHEN OTHERS =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001");
        state_var_NS <= for_C_0;
    END CASE;
  END PROCESS fir_core_core_fsm_1;

  fir_core_core_fsm_1_REG : PROCESS (clk)
  BEGIN
    IF clk'event AND ( clk = '1' ) THEN
      IF ( rst = '1' ) THEN
        state_var <= main_C_0;
      ELSE
        state_var <= state_var_NS;
      END IF;
    END IF;
  END PROCESS fir_core_core_fsm_1_REG;

END v1;

-- ------------------------------------------------------------------
--  Design Unit:    fir_core
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.ccs_out_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;


ENTITY fir_core IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    input_rsc_dat : IN STD_LOGIC_VECTOR (4095 DOWNTO 0);
    input_rsc_triosy_lz : OUT STD_LOGIC;
    output_rsc_dat : OUT STD_LOGIC_VECTOR (4095 DOWNTO 0);
    output_rsc_triosy_lz : OUT STD_LOGIC
  );
END fir_core;

ARCHITECTURE v1 OF fir_core IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL input_rsci_idat : STD_LOGIC_VECTOR (4095 DOWNTO 0);
  SIGNAL output_rsci_idat_4095_4064 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_4063_4032 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_4031_4000 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_3999_3968 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_3967_3936 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_3935_3904 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_3903_3872 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_3871_3840 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_3839_3808 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_3807_3776 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_3775_3744 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_3743_3712 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_3711_3680 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_3679_3648 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_3647_3616 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_3615_3584 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_3583_3552 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_3551_3520 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_3519_3488 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_3487_3456 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_3455_3424 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_3423_3392 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_3391_3360 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_3359_3328 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_3327_3296 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_3295_3264 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_3263_3232 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_3231_3200 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_3199_3168 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_3167_3136 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_3135_3104 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_3103_3072 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_3071_3040 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_3039_3008 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_3007_2976 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_2975_2944 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_2943_2912 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_2911_2880 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_2879_2848 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_2847_2816 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_2815_2784 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_2783_2752 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_2751_2720 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_2719_2688 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_2687_2656 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_2655_2624 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_2623_2592 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_2591_2560 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_2559_2528 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_2527_2496 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_2495_2464 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_2463_2432 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_2431_2400 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_2399_2368 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_2367_2336 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_2335_2304 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_2303_2272 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_2271_2240 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_2239_2208 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_2207_2176 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_2175_2144 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_2143_2112 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_2111_2080 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_2079_2048 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_2047_2016 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_2015_1984 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_1983_1952 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_1951_1920 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_1919_1888 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_1887_1856 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_1855_1824 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_1823_1792 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_1791_1760 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_1759_1728 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_1727_1696 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_1695_1664 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_1663_1632 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_1631_1600 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_1599_1568 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_1567_1536 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_1535_1504 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_1503_1472 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_1471_1440 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_1439_1408 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_1407_1376 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_1375_1344 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_1343_1312 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_1311_1280 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_1279_1248 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_1247_1216 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_1215_1184 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_1183_1152 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_1151_1120 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_1119_1088 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_1087_1056 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_1055_1024 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_1023_992 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_991_960 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_959_928 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_927_896 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_895_864 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_863_832 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_831_800 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_799_768 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_767_736 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_735_704 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_703_672 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_671_640 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_639_608 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_607_576 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_575_544 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_543_512 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_511_480 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_479_448 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_447_416 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_415_384 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_383_352 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_351_320 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_319_288 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_287_256 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_255_224 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_223_192 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_191_160 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_159_128 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_127_96 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_95_64 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_63_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsci_idat_31_0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL fsm_output : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL for_or_tmp : STD_LOGIC;
  SIGNAL or_dcpl_330 : STD_LOGIC;
  SIGNAL or_dcpl_331 : STD_LOGIC;
  SIGNAL or_dcpl_332 : STD_LOGIC;
  SIGNAL or_dcpl_333 : STD_LOGIC;
  SIGNAL or_dcpl_334 : STD_LOGIC;
  SIGNAL or_dcpl_335 : STD_LOGIC;
  SIGNAL or_dcpl_336 : STD_LOGIC;
  SIGNAL or_tmp_259 : STD_LOGIC;
  SIGNAL or_tmp_643 : STD_LOGIC;
  SIGNAL for_nor_62_itm : STD_LOGIC;
  SIGNAL for_nor_31_itm : STD_LOGIC;
  SIGNAL for_nor_15_itm : STD_LOGIC;
  SIGNAL for_nor_7_itm : STD_LOGIC;
  SIGNAL for_nor_3_itm : STD_LOGIC;
  SIGNAL for_nor_1_itm : STD_LOGIC;
  SIGNAL for_nor_itm : STD_LOGIC;
  SIGNAL i_7_0_sva_6_0 : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL i_7_0_sva_1 : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL for_equal_tmp_3 : STD_LOGIC;
  SIGNAL for_equal_tmp_5 : STD_LOGIC;
  SIGNAL for_equal_tmp_6 : STD_LOGIC;
  SIGNAL for_equal_tmp_7 : STD_LOGIC;
  SIGNAL for_equal_tmp_9 : STD_LOGIC;
  SIGNAL for_equal_tmp_10 : STD_LOGIC;
  SIGNAL for_equal_tmp_11 : STD_LOGIC;
  SIGNAL for_equal_tmp_12 : STD_LOGIC;
  SIGNAL for_equal_tmp_13 : STD_LOGIC;
  SIGNAL for_equal_tmp_14 : STD_LOGIC;
  SIGNAL for_equal_tmp_15 : STD_LOGIC;
  SIGNAL for_equal_tmp_17 : STD_LOGIC;
  SIGNAL for_equal_tmp_18 : STD_LOGIC;
  SIGNAL for_equal_tmp_19 : STD_LOGIC;
  SIGNAL for_equal_tmp_20 : STD_LOGIC;
  SIGNAL for_equal_tmp_21 : STD_LOGIC;
  SIGNAL for_equal_tmp_22 : STD_LOGIC;
  SIGNAL for_equal_tmp_23 : STD_LOGIC;
  SIGNAL for_equal_tmp_24 : STD_LOGIC;
  SIGNAL for_equal_tmp_25 : STD_LOGIC;
  SIGNAL for_equal_tmp_26 : STD_LOGIC;
  SIGNAL for_equal_tmp_27 : STD_LOGIC;
  SIGNAL for_equal_tmp_28 : STD_LOGIC;
  SIGNAL for_equal_tmp_29 : STD_LOGIC;
  SIGNAL for_equal_tmp_30 : STD_LOGIC;
  SIGNAL for_equal_tmp_31 : STD_LOGIC;
  SIGNAL for_equal_tmp_33 : STD_LOGIC;
  SIGNAL for_equal_tmp_34 : STD_LOGIC;
  SIGNAL for_equal_tmp_35 : STD_LOGIC;
  SIGNAL for_equal_tmp_36 : STD_LOGIC;
  SIGNAL for_equal_tmp_37 : STD_LOGIC;
  SIGNAL for_equal_tmp_38 : STD_LOGIC;
  SIGNAL for_equal_tmp_39 : STD_LOGIC;
  SIGNAL for_equal_tmp_40 : STD_LOGIC;
  SIGNAL for_equal_tmp_41 : STD_LOGIC;
  SIGNAL for_equal_tmp_42 : STD_LOGIC;
  SIGNAL for_equal_tmp_43 : STD_LOGIC;
  SIGNAL for_equal_tmp_44 : STD_LOGIC;
  SIGNAL for_equal_tmp_45 : STD_LOGIC;
  SIGNAL for_equal_tmp_46 : STD_LOGIC;
  SIGNAL for_equal_tmp_47 : STD_LOGIC;
  SIGNAL for_equal_tmp_48 : STD_LOGIC;
  SIGNAL for_equal_tmp_49 : STD_LOGIC;
  SIGNAL for_equal_tmp_50 : STD_LOGIC;
  SIGNAL for_equal_tmp_51 : STD_LOGIC;
  SIGNAL for_equal_tmp_52 : STD_LOGIC;
  SIGNAL for_equal_tmp_53 : STD_LOGIC;
  SIGNAL for_equal_tmp_54 : STD_LOGIC;
  SIGNAL for_equal_tmp_55 : STD_LOGIC;
  SIGNAL for_equal_tmp_56 : STD_LOGIC;
  SIGNAL for_equal_tmp_57 : STD_LOGIC;
  SIGNAL for_equal_tmp_58 : STD_LOGIC;
  SIGNAL for_equal_tmp_59 : STD_LOGIC;
  SIGNAL for_equal_tmp_60 : STD_LOGIC;
  SIGNAL for_equal_tmp_61 : STD_LOGIC;
  SIGNAL for_equal_tmp_62 : STD_LOGIC;
  SIGNAL for_equal_tmp_63 : STD_LOGIC;
  SIGNAL for_equal_tmp_65 : STD_LOGIC;
  SIGNAL for_equal_tmp_66 : STD_LOGIC;
  SIGNAL for_equal_tmp_67 : STD_LOGIC;
  SIGNAL for_equal_tmp_68 : STD_LOGIC;
  SIGNAL for_equal_tmp_69 : STD_LOGIC;
  SIGNAL for_equal_tmp_70 : STD_LOGIC;
  SIGNAL for_equal_tmp_71 : STD_LOGIC;
  SIGNAL for_equal_tmp_72 : STD_LOGIC;
  SIGNAL for_equal_tmp_73 : STD_LOGIC;
  SIGNAL for_equal_tmp_74 : STD_LOGIC;
  SIGNAL for_equal_tmp_75 : STD_LOGIC;
  SIGNAL for_equal_tmp_76 : STD_LOGIC;
  SIGNAL for_equal_tmp_77 : STD_LOGIC;
  SIGNAL for_equal_tmp_78 : STD_LOGIC;
  SIGNAL for_equal_tmp_79 : STD_LOGIC;
  SIGNAL for_equal_tmp_80 : STD_LOGIC;
  SIGNAL for_equal_tmp_81 : STD_LOGIC;
  SIGNAL for_equal_tmp_82 : STD_LOGIC;
  SIGNAL for_equal_tmp_83 : STD_LOGIC;
  SIGNAL for_equal_tmp_84 : STD_LOGIC;
  SIGNAL for_equal_tmp_85 : STD_LOGIC;
  SIGNAL for_equal_tmp_86 : STD_LOGIC;
  SIGNAL for_equal_tmp_87 : STD_LOGIC;
  SIGNAL for_equal_tmp_88 : STD_LOGIC;
  SIGNAL for_equal_tmp_89 : STD_LOGIC;
  SIGNAL for_equal_tmp_90 : STD_LOGIC;
  SIGNAL for_equal_tmp_91 : STD_LOGIC;
  SIGNAL for_equal_tmp_92 : STD_LOGIC;
  SIGNAL for_equal_tmp_93 : STD_LOGIC;
  SIGNAL for_equal_tmp_94 : STD_LOGIC;
  SIGNAL for_equal_tmp_95 : STD_LOGIC;
  SIGNAL for_equal_tmp_96 : STD_LOGIC;
  SIGNAL for_equal_tmp_97 : STD_LOGIC;
  SIGNAL for_equal_tmp_98 : STD_LOGIC;
  SIGNAL for_equal_tmp_99 : STD_LOGIC;
  SIGNAL for_equal_tmp_100 : STD_LOGIC;
  SIGNAL for_equal_tmp_101 : STD_LOGIC;
  SIGNAL for_equal_tmp_102 : STD_LOGIC;
  SIGNAL for_equal_tmp_103 : STD_LOGIC;
  SIGNAL for_equal_tmp_104 : STD_LOGIC;
  SIGNAL for_equal_tmp_105 : STD_LOGIC;
  SIGNAL for_equal_tmp_106 : STD_LOGIC;
  SIGNAL for_equal_tmp_107 : STD_LOGIC;
  SIGNAL for_equal_tmp_108 : STD_LOGIC;
  SIGNAL for_equal_tmp_109 : STD_LOGIC;
  SIGNAL for_equal_tmp_110 : STD_LOGIC;
  SIGNAL for_equal_tmp_111 : STD_LOGIC;
  SIGNAL for_equal_tmp_112 : STD_LOGIC;
  SIGNAL for_equal_tmp_113 : STD_LOGIC;
  SIGNAL for_equal_tmp_114 : STD_LOGIC;
  SIGNAL for_equal_tmp_115 : STD_LOGIC;
  SIGNAL for_equal_tmp_116 : STD_LOGIC;
  SIGNAL for_equal_tmp_117 : STD_LOGIC;
  SIGNAL for_equal_tmp_118 : STD_LOGIC;
  SIGNAL for_equal_tmp_119 : STD_LOGIC;
  SIGNAL for_equal_tmp_120 : STD_LOGIC;
  SIGNAL for_equal_tmp_121 : STD_LOGIC;
  SIGNAL for_equal_tmp_122 : STD_LOGIC;
  SIGNAL for_equal_tmp_123 : STD_LOGIC;
  SIGNAL for_equal_tmp_124 : STD_LOGIC;
  SIGNAL for_equal_tmp_125 : STD_LOGIC;
  SIGNAL for_equal_tmp_126 : STD_LOGIC;
  SIGNAL for_equal_tmp_127 : STD_LOGIC;
  SIGNAL reg_output_rsc_triosy_obj_ld_cse : STD_LOGIC;
  SIGNAL output_output_mux_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_2047_2016_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_2079_2048_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_2015_1984_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_2111_2080_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_1983_1952_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_2143_2112_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_1951_1920_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_2175_2144_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_1919_1888_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_2207_2176_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_1887_1856_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_2239_2208_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_1855_1824_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_2271_2240_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_1823_1792_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_2303_2272_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_1791_1760_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_2335_2304_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_1759_1728_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_2367_2336_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_1727_1696_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_2399_2368_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_1695_1664_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_2431_2400_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_1663_1632_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_2463_2432_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_1631_1600_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_2495_2464_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_1599_1568_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_2527_2496_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_1567_1536_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_2559_2528_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_1535_1504_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_2591_2560_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_1503_1472_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_2623_2592_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_1471_1440_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_2655_2624_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_1439_1408_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_2687_2656_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_1407_1376_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_2719_2688_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_1375_1344_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_2751_2720_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_1343_1312_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_2783_2752_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_1311_1280_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_2815_2784_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_1279_1248_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_2847_2816_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_1247_1216_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_2879_2848_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_1215_1184_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_2911_2880_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_1183_1152_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_2943_2912_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_1151_1120_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_2975_2944_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_1119_1088_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_3007_2976_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_1087_1056_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_3039_3008_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_1055_1024_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_3071_3040_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_1023_992_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_3103_3072_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_991_960_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_3135_3104_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_959_928_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_3167_3136_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_927_896_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_3199_3168_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_895_864_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_3231_3200_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_863_832_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_3263_3232_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_831_800_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_3295_3264_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_799_768_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_3327_3296_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_767_736_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_3359_3328_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_735_704_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_3391_3360_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_703_672_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_3423_3392_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_671_640_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_3455_3424_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_639_608_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_3487_3456_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_607_576_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_3519_3488_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_575_544_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_3551_3520_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_543_512_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_3583_3552_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_511_480_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_3615_3584_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_479_448_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_3647_3616_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_447_416_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_3679_3648_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_415_384_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_3711_3680_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_383_352_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_3743_3712_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_351_320_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_3775_3744_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_319_288_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_3807_3776_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_287_256_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_3839_3808_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_255_224_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_3871_3840_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_223_192_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_3903_3872_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_191_160_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_3935_3904_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_159_128_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_3967_3936_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_127_96_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_3999_3968_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_95_64_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_4031_4000_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_63_32_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_4063_4032_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_31_0_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL output_rsc_1_4095_4064_lpi_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL for_io_read_output_rsc_sdt_4095_4064_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_4063_4032_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_4031_4000_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_3999_3968_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_3967_3936_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_3935_3904_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_3903_3872_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_3871_3840_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_3839_3808_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_3807_3776_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_3775_3744_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_3743_3712_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_3711_3680_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_3679_3648_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_3647_3616_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_3615_3584_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_3583_3552_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_3551_3520_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_3519_3488_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_3487_3456_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_3455_3424_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_3423_3392_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_3391_3360_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_3359_3328_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_3327_3296_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_3295_3264_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_3263_3232_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_3231_3200_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_3199_3168_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_3167_3136_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_3135_3104_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_3103_3072_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_3071_3040_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_3039_3008_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_3007_2976_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_2975_2944_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_2943_2912_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_2911_2880_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_2879_2848_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_2847_2816_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_2815_2784_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_2783_2752_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_2751_2720_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_2719_2688_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_2687_2656_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_2655_2624_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_2623_2592_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_2591_2560_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_2559_2528_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_2527_2496_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_2495_2464_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_2463_2432_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_2431_2400_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_2399_2368_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_2367_2336_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_2335_2304_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_2303_2272_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_2271_2240_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_2239_2208_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_2207_2176_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_2175_2144_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_2143_2112_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_2111_2080_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_2079_2048_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_2047_2016_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_2015_1984_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_1983_1952_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_1951_1920_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_1919_1888_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_1887_1856_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_1855_1824_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_1823_1792_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_1791_1760_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_1759_1728_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_1727_1696_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_1695_1664_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_1663_1632_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_1631_1600_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_1599_1568_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_1567_1536_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_1535_1504_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_1503_1472_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_1471_1440_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_1439_1408_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_1407_1376_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_1375_1344_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_1343_1312_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_1311_1280_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_1279_1248_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_1247_1216_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_1215_1184_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_1183_1152_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_1151_1120_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_1119_1088_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_1087_1056_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_1055_1024_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_1023_992_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_991_960_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_959_928_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_927_896_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_895_864_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_863_832_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_831_800_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_799_768_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_767_736_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_735_704_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_703_672_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_671_640_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_639_608_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_607_576_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_575_544_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_543_512_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_511_480_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_479_448_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_447_416_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_415_384_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_383_352_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_351_320_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_319_288_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_287_256_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_255_224_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_223_192_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_191_160_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_159_128_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_127_96_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_95_64_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_63_32_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_io_read_output_rsc_sdt_31_0_lpi_2_dfm : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL for_mux_itm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL for_for_mul_1_cmx_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_output_rsc_1_31_output_or_cse : STD_LOGIC;

  SIGNAL and_660_nl : STD_LOGIC;
  SIGNAL and_666_nl : STD_LOGIC;
  SIGNAL and_672_nl : STD_LOGIC;
  SIGNAL and_678_nl : STD_LOGIC;
  SIGNAL and_684_nl : STD_LOGIC;
  SIGNAL and_690_nl : STD_LOGIC;
  SIGNAL and_696_nl : STD_LOGIC;
  SIGNAL and_702_nl : STD_LOGIC;
  SIGNAL and_708_nl : STD_LOGIC;
  SIGNAL and_714_nl : STD_LOGIC;
  SIGNAL and_720_nl : STD_LOGIC;
  SIGNAL and_726_nl : STD_LOGIC;
  SIGNAL and_732_nl : STD_LOGIC;
  SIGNAL and_738_nl : STD_LOGIC;
  SIGNAL and_744_nl : STD_LOGIC;
  SIGNAL and_750_nl : STD_LOGIC;
  SIGNAL and_756_nl : STD_LOGIC;
  SIGNAL and_762_nl : STD_LOGIC;
  SIGNAL and_768_nl : STD_LOGIC;
  SIGNAL and_774_nl : STD_LOGIC;
  SIGNAL and_780_nl : STD_LOGIC;
  SIGNAL and_786_nl : STD_LOGIC;
  SIGNAL and_792_nl : STD_LOGIC;
  SIGNAL and_798_nl : STD_LOGIC;
  SIGNAL and_804_nl : STD_LOGIC;
  SIGNAL and_810_nl : STD_LOGIC;
  SIGNAL and_816_nl : STD_LOGIC;
  SIGNAL and_822_nl : STD_LOGIC;
  SIGNAL and_828_nl : STD_LOGIC;
  SIGNAL and_834_nl : STD_LOGIC;
  SIGNAL and_840_nl : STD_LOGIC;
  SIGNAL and_846_nl : STD_LOGIC;
  SIGNAL and_852_nl : STD_LOGIC;
  SIGNAL and_858_nl : STD_LOGIC;
  SIGNAL and_864_nl : STD_LOGIC;
  SIGNAL and_870_nl : STD_LOGIC;
  SIGNAL and_876_nl : STD_LOGIC;
  SIGNAL and_882_nl : STD_LOGIC;
  SIGNAL and_888_nl : STD_LOGIC;
  SIGNAL and_894_nl : STD_LOGIC;
  SIGNAL and_900_nl : STD_LOGIC;
  SIGNAL and_906_nl : STD_LOGIC;
  SIGNAL and_912_nl : STD_LOGIC;
  SIGNAL and_918_nl : STD_LOGIC;
  SIGNAL and_924_nl : STD_LOGIC;
  SIGNAL and_930_nl : STD_LOGIC;
  SIGNAL and_936_nl : STD_LOGIC;
  SIGNAL and_942_nl : STD_LOGIC;
  SIGNAL and_948_nl : STD_LOGIC;
  SIGNAL and_954_nl : STD_LOGIC;
  SIGNAL and_960_nl : STD_LOGIC;
  SIGNAL and_966_nl : STD_LOGIC;
  SIGNAL and_972_nl : STD_LOGIC;
  SIGNAL and_978_nl : STD_LOGIC;
  SIGNAL and_984_nl : STD_LOGIC;
  SIGNAL and_990_nl : STD_LOGIC;
  SIGNAL and_996_nl : STD_LOGIC;
  SIGNAL and_1002_nl : STD_LOGIC;
  SIGNAL and_1008_nl : STD_LOGIC;
  SIGNAL and_1014_nl : STD_LOGIC;
  SIGNAL and_1020_nl : STD_LOGIC;
  SIGNAL and_1026_nl : STD_LOGIC;
  SIGNAL and_1032_nl : STD_LOGIC;
  SIGNAL and_1038_nl : STD_LOGIC;
  SIGNAL and_1044_nl : STD_LOGIC;
  SIGNAL and_1050_nl : STD_LOGIC;
  SIGNAL and_1056_nl : STD_LOGIC;
  SIGNAL and_1062_nl : STD_LOGIC;
  SIGNAL and_1068_nl : STD_LOGIC;
  SIGNAL and_1074_nl : STD_LOGIC;
  SIGNAL and_1080_nl : STD_LOGIC;
  SIGNAL and_1086_nl : STD_LOGIC;
  SIGNAL and_1092_nl : STD_LOGIC;
  SIGNAL and_1098_nl : STD_LOGIC;
  SIGNAL and_1104_nl : STD_LOGIC;
  SIGNAL and_1110_nl : STD_LOGIC;
  SIGNAL and_1116_nl : STD_LOGIC;
  SIGNAL and_1122_nl : STD_LOGIC;
  SIGNAL and_1128_nl : STD_LOGIC;
  SIGNAL and_1134_nl : STD_LOGIC;
  SIGNAL and_1140_nl : STD_LOGIC;
  SIGNAL and_1146_nl : STD_LOGIC;
  SIGNAL and_1152_nl : STD_LOGIC;
  SIGNAL and_1158_nl : STD_LOGIC;
  SIGNAL and_1164_nl : STD_LOGIC;
  SIGNAL and_1170_nl : STD_LOGIC;
  SIGNAL and_1176_nl : STD_LOGIC;
  SIGNAL and_1182_nl : STD_LOGIC;
  SIGNAL and_1188_nl : STD_LOGIC;
  SIGNAL and_1194_nl : STD_LOGIC;
  SIGNAL and_1200_nl : STD_LOGIC;
  SIGNAL and_1206_nl : STD_LOGIC;
  SIGNAL and_1212_nl : STD_LOGIC;
  SIGNAL and_1218_nl : STD_LOGIC;
  SIGNAL and_1224_nl : STD_LOGIC;
  SIGNAL and_1230_nl : STD_LOGIC;
  SIGNAL and_1236_nl : STD_LOGIC;
  SIGNAL and_1242_nl : STD_LOGIC;
  SIGNAL and_1248_nl : STD_LOGIC;
  SIGNAL and_1254_nl : STD_LOGIC;
  SIGNAL and_1260_nl : STD_LOGIC;
  SIGNAL and_1266_nl : STD_LOGIC;
  SIGNAL and_1272_nl : STD_LOGIC;
  SIGNAL and_1278_nl : STD_LOGIC;
  SIGNAL and_1284_nl : STD_LOGIC;
  SIGNAL and_1290_nl : STD_LOGIC;
  SIGNAL and_1296_nl : STD_LOGIC;
  SIGNAL and_1302_nl : STD_LOGIC;
  SIGNAL and_1308_nl : STD_LOGIC;
  SIGNAL and_1314_nl : STD_LOGIC;
  SIGNAL and_1320_nl : STD_LOGIC;
  SIGNAL and_1326_nl : STD_LOGIC;
  SIGNAL and_1332_nl : STD_LOGIC;
  SIGNAL and_1338_nl : STD_LOGIC;
  SIGNAL and_1344_nl : STD_LOGIC;
  SIGNAL and_1350_nl : STD_LOGIC;
  SIGNAL and_1356_nl : STD_LOGIC;
  SIGNAL and_1362_nl : STD_LOGIC;
  SIGNAL and_1368_nl : STD_LOGIC;
  SIGNAL and_1374_nl : STD_LOGIC;
  SIGNAL and_1380_nl : STD_LOGIC;
  SIGNAL and_1386_nl : STD_LOGIC;
  SIGNAL and_1392_nl : STD_LOGIC;
  SIGNAL and_1398_nl : STD_LOGIC;
  SIGNAL and_1404_nl : STD_LOGIC;
  SIGNAL and_1410_nl : STD_LOGIC;
  SIGNAL and_1416_nl : STD_LOGIC;
  SIGNAL for_and_253_nl : STD_LOGIC;
  SIGNAL for_and_251_nl : STD_LOGIC;
  SIGNAL for_and_249_nl : STD_LOGIC;
  SIGNAL for_and_247_nl : STD_LOGIC;
  SIGNAL for_and_245_nl : STD_LOGIC;
  SIGNAL for_and_243_nl : STD_LOGIC;
  SIGNAL for_and_241_nl : STD_LOGIC;
  SIGNAL for_and_239_nl : STD_LOGIC;
  SIGNAL for_and_237_nl : STD_LOGIC;
  SIGNAL for_and_235_nl : STD_LOGIC;
  SIGNAL for_and_233_nl : STD_LOGIC;
  SIGNAL for_and_231_nl : STD_LOGIC;
  SIGNAL for_and_229_nl : STD_LOGIC;
  SIGNAL for_and_227_nl : STD_LOGIC;
  SIGNAL for_and_225_nl : STD_LOGIC;
  SIGNAL for_and_223_nl : STD_LOGIC;
  SIGNAL for_and_221_nl : STD_LOGIC;
  SIGNAL for_and_219_nl : STD_LOGIC;
  SIGNAL for_and_217_nl : STD_LOGIC;
  SIGNAL for_and_215_nl : STD_LOGIC;
  SIGNAL for_and_213_nl : STD_LOGIC;
  SIGNAL for_and_211_nl : STD_LOGIC;
  SIGNAL for_and_209_nl : STD_LOGIC;
  SIGNAL for_and_207_nl : STD_LOGIC;
  SIGNAL for_and_205_nl : STD_LOGIC;
  SIGNAL for_and_203_nl : STD_LOGIC;
  SIGNAL for_and_201_nl : STD_LOGIC;
  SIGNAL for_and_199_nl : STD_LOGIC;
  SIGNAL for_and_197_nl : STD_LOGIC;
  SIGNAL for_and_195_nl : STD_LOGIC;
  SIGNAL for_and_193_nl : STD_LOGIC;
  SIGNAL for_and_191_nl : STD_LOGIC;
  SIGNAL for_and_189_nl : STD_LOGIC;
  SIGNAL for_and_187_nl : STD_LOGIC;
  SIGNAL for_and_185_nl : STD_LOGIC;
  SIGNAL for_and_183_nl : STD_LOGIC;
  SIGNAL for_and_181_nl : STD_LOGIC;
  SIGNAL for_and_179_nl : STD_LOGIC;
  SIGNAL for_and_177_nl : STD_LOGIC;
  SIGNAL for_and_175_nl : STD_LOGIC;
  SIGNAL for_and_173_nl : STD_LOGIC;
  SIGNAL for_and_171_nl : STD_LOGIC;
  SIGNAL for_and_169_nl : STD_LOGIC;
  SIGNAL for_and_167_nl : STD_LOGIC;
  SIGNAL for_and_165_nl : STD_LOGIC;
  SIGNAL for_and_163_nl : STD_LOGIC;
  SIGNAL for_and_161_nl : STD_LOGIC;
  SIGNAL for_and_159_nl : STD_LOGIC;
  SIGNAL for_and_157_nl : STD_LOGIC;
  SIGNAL for_and_155_nl : STD_LOGIC;
  SIGNAL for_and_153_nl : STD_LOGIC;
  SIGNAL for_and_151_nl : STD_LOGIC;
  SIGNAL for_and_149_nl : STD_LOGIC;
  SIGNAL for_and_147_nl : STD_LOGIC;
  SIGNAL for_and_145_nl : STD_LOGIC;
  SIGNAL for_and_143_nl : STD_LOGIC;
  SIGNAL for_and_141_nl : STD_LOGIC;
  SIGNAL for_and_139_nl : STD_LOGIC;
  SIGNAL for_and_137_nl : STD_LOGIC;
  SIGNAL for_and_135_nl : STD_LOGIC;
  SIGNAL for_and_133_nl : STD_LOGIC;
  SIGNAL for_and_131_nl : STD_LOGIC;
  SIGNAL for_and_129_nl : STD_LOGIC;
  SIGNAL for_and_127_nl : STD_LOGIC;
  SIGNAL for_and_125_nl : STD_LOGIC;
  SIGNAL for_and_123_nl : STD_LOGIC;
  SIGNAL for_and_121_nl : STD_LOGIC;
  SIGNAL for_and_119_nl : STD_LOGIC;
  SIGNAL for_and_117_nl : STD_LOGIC;
  SIGNAL for_and_115_nl : STD_LOGIC;
  SIGNAL for_and_113_nl : STD_LOGIC;
  SIGNAL for_and_111_nl : STD_LOGIC;
  SIGNAL for_and_109_nl : STD_LOGIC;
  SIGNAL for_and_107_nl : STD_LOGIC;
  SIGNAL for_and_105_nl : STD_LOGIC;
  SIGNAL for_and_103_nl : STD_LOGIC;
  SIGNAL for_and_101_nl : STD_LOGIC;
  SIGNAL for_and_99_nl : STD_LOGIC;
  SIGNAL for_and_97_nl : STD_LOGIC;
  SIGNAL for_and_95_nl : STD_LOGIC;
  SIGNAL for_and_93_nl : STD_LOGIC;
  SIGNAL for_and_91_nl : STD_LOGIC;
  SIGNAL for_and_89_nl : STD_LOGIC;
  SIGNAL for_and_87_nl : STD_LOGIC;
  SIGNAL for_and_85_nl : STD_LOGIC;
  SIGNAL for_and_83_nl : STD_LOGIC;
  SIGNAL for_and_81_nl : STD_LOGIC;
  SIGNAL for_and_79_nl : STD_LOGIC;
  SIGNAL for_and_77_nl : STD_LOGIC;
  SIGNAL for_and_75_nl : STD_LOGIC;
  SIGNAL for_and_73_nl : STD_LOGIC;
  SIGNAL for_and_71_nl : STD_LOGIC;
  SIGNAL for_and_69_nl : STD_LOGIC;
  SIGNAL for_and_67_nl : STD_LOGIC;
  SIGNAL for_and_65_nl : STD_LOGIC;
  SIGNAL for_and_63_nl : STD_LOGIC;
  SIGNAL for_and_61_nl : STD_LOGIC;
  SIGNAL for_and_59_nl : STD_LOGIC;
  SIGNAL for_and_57_nl : STD_LOGIC;
  SIGNAL for_and_55_nl : STD_LOGIC;
  SIGNAL for_and_53_nl : STD_LOGIC;
  SIGNAL for_and_51_nl : STD_LOGIC;
  SIGNAL for_and_49_nl : STD_LOGIC;
  SIGNAL for_and_47_nl : STD_LOGIC;
  SIGNAL for_and_45_nl : STD_LOGIC;
  SIGNAL for_and_43_nl : STD_LOGIC;
  SIGNAL for_and_41_nl : STD_LOGIC;
  SIGNAL for_and_39_nl : STD_LOGIC;
  SIGNAL for_and_37_nl : STD_LOGIC;
  SIGNAL for_and_35_nl : STD_LOGIC;
  SIGNAL for_and_33_nl : STD_LOGIC;
  SIGNAL for_and_31_nl : STD_LOGIC;
  SIGNAL for_and_29_nl : STD_LOGIC;
  SIGNAL for_and_27_nl : STD_LOGIC;
  SIGNAL for_and_25_nl : STD_LOGIC;
  SIGNAL for_and_23_nl : STD_LOGIC;
  SIGNAL for_and_21_nl : STD_LOGIC;
  SIGNAL for_and_19_nl : STD_LOGIC;
  SIGNAL for_and_17_nl : STD_LOGIC;
  SIGNAL for_and_15_nl : STD_LOGIC;
  SIGNAL for_and_13_nl : STD_LOGIC;
  SIGNAL for_and_11_nl : STD_LOGIC;
  SIGNAL for_and_9_nl : STD_LOGIC;
  SIGNAL for_and_7_nl : STD_LOGIC;
  SIGNAL for_and_5_nl : STD_LOGIC;
  SIGNAL for_and_3_nl : STD_LOGIC;
  SIGNAL for_and_1_nl : STD_LOGIC;
  SIGNAL input_rsci_dat : STD_LOGIC_VECTOR (4095 DOWNTO 0);
  SIGNAL input_rsci_idat_1 : STD_LOGIC_VECTOR (4095 DOWNTO 0);

  SIGNAL output_rsci_idat : STD_LOGIC_VECTOR (4095 DOWNTO 0);
  SIGNAL output_rsci_dat : STD_LOGIC_VECTOR (4095 DOWNTO 0);

  COMPONENT fir_core_core_fsm
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      fsm_output : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      for_C_2_tr0 : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL fir_core_core_fsm_inst_fsm_output : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL fir_core_core_fsm_inst_for_C_2_tr0 : STD_LOGIC;

  FUNCTION CONV_SL_1_1(input_val:BOOLEAN)
  RETURN STD_LOGIC IS
  BEGIN
    IF input_val THEN RETURN '1';ELSE RETURN '0';END IF;
  END;

  FUNCTION MUX_v_32_128_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_15 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_16 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_17 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_18 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_19 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_20 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_21 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_22 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_23 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_24 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_25 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_26 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_27 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_28 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_29 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_30 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_31 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_32 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_33 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_34 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_35 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_36 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_37 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_38 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_39 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_40 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_41 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_42 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_43 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_44 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_45 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_46 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_47 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_48 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_49 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_50 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_51 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_52 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_53 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_54 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_55 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_56 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_57 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_58 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_59 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_60 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_61 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_62 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_63 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_64 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_65 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_66 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_67 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_68 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_69 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_70 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_71 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_72 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_73 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_74 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_75 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_76 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_77 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_78 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_79 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_80 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_81 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_82 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_83 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_84 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_85 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_86 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_87 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_88 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_89 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_90 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_91 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_92 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_93 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_94 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_95 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_96 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_97 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_98 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_99 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_100 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_101 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_102 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_103 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_104 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_105 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_106 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_107 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_108 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_109 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_110 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_111 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_112 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_113 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_114 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_115 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_116 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_117 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_118 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_119 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_120 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_121 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_122 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_123 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_124 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_125 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_126 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_127 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(6 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN "0000000" =>
          result := input_0;
        WHEN "0000001" =>
          result := input_1;
        WHEN "0000010" =>
          result := input_2;
        WHEN "0000011" =>
          result := input_3;
        WHEN "0000100" =>
          result := input_4;
        WHEN "0000101" =>
          result := input_5;
        WHEN "0000110" =>
          result := input_6;
        WHEN "0000111" =>
          result := input_7;
        WHEN "0001000" =>
          result := input_8;
        WHEN "0001001" =>
          result := input_9;
        WHEN "0001010" =>
          result := input_10;
        WHEN "0001011" =>
          result := input_11;
        WHEN "0001100" =>
          result := input_12;
        WHEN "0001101" =>
          result := input_13;
        WHEN "0001110" =>
          result := input_14;
        WHEN "0001111" =>
          result := input_15;
        WHEN "0010000" =>
          result := input_16;
        WHEN "0010001" =>
          result := input_17;
        WHEN "0010010" =>
          result := input_18;
        WHEN "0010011" =>
          result := input_19;
        WHEN "0010100" =>
          result := input_20;
        WHEN "0010101" =>
          result := input_21;
        WHEN "0010110" =>
          result := input_22;
        WHEN "0010111" =>
          result := input_23;
        WHEN "0011000" =>
          result := input_24;
        WHEN "0011001" =>
          result := input_25;
        WHEN "0011010" =>
          result := input_26;
        WHEN "0011011" =>
          result := input_27;
        WHEN "0011100" =>
          result := input_28;
        WHEN "0011101" =>
          result := input_29;
        WHEN "0011110" =>
          result := input_30;
        WHEN "0011111" =>
          result := input_31;
        WHEN "0100000" =>
          result := input_32;
        WHEN "0100001" =>
          result := input_33;
        WHEN "0100010" =>
          result := input_34;
        WHEN "0100011" =>
          result := input_35;
        WHEN "0100100" =>
          result := input_36;
        WHEN "0100101" =>
          result := input_37;
        WHEN "0100110" =>
          result := input_38;
        WHEN "0100111" =>
          result := input_39;
        WHEN "0101000" =>
          result := input_40;
        WHEN "0101001" =>
          result := input_41;
        WHEN "0101010" =>
          result := input_42;
        WHEN "0101011" =>
          result := input_43;
        WHEN "0101100" =>
          result := input_44;
        WHEN "0101101" =>
          result := input_45;
        WHEN "0101110" =>
          result := input_46;
        WHEN "0101111" =>
          result := input_47;
        WHEN "0110000" =>
          result := input_48;
        WHEN "0110001" =>
          result := input_49;
        WHEN "0110010" =>
          result := input_50;
        WHEN "0110011" =>
          result := input_51;
        WHEN "0110100" =>
          result := input_52;
        WHEN "0110101" =>
          result := input_53;
        WHEN "0110110" =>
          result := input_54;
        WHEN "0110111" =>
          result := input_55;
        WHEN "0111000" =>
          result := input_56;
        WHEN "0111001" =>
          result := input_57;
        WHEN "0111010" =>
          result := input_58;
        WHEN "0111011" =>
          result := input_59;
        WHEN "0111100" =>
          result := input_60;
        WHEN "0111101" =>
          result := input_61;
        WHEN "0111110" =>
          result := input_62;
        WHEN "0111111" =>
          result := input_63;
        WHEN "1000000" =>
          result := input_64;
        WHEN "1000001" =>
          result := input_65;
        WHEN "1000010" =>
          result := input_66;
        WHEN "1000011" =>
          result := input_67;
        WHEN "1000100" =>
          result := input_68;
        WHEN "1000101" =>
          result := input_69;
        WHEN "1000110" =>
          result := input_70;
        WHEN "1000111" =>
          result := input_71;
        WHEN "1001000" =>
          result := input_72;
        WHEN "1001001" =>
          result := input_73;
        WHEN "1001010" =>
          result := input_74;
        WHEN "1001011" =>
          result := input_75;
        WHEN "1001100" =>
          result := input_76;
        WHEN "1001101" =>
          result := input_77;
        WHEN "1001110" =>
          result := input_78;
        WHEN "1001111" =>
          result := input_79;
        WHEN "1010000" =>
          result := input_80;
        WHEN "1010001" =>
          result := input_81;
        WHEN "1010010" =>
          result := input_82;
        WHEN "1010011" =>
          result := input_83;
        WHEN "1010100" =>
          result := input_84;
        WHEN "1010101" =>
          result := input_85;
        WHEN "1010110" =>
          result := input_86;
        WHEN "1010111" =>
          result := input_87;
        WHEN "1011000" =>
          result := input_88;
        WHEN "1011001" =>
          result := input_89;
        WHEN "1011010" =>
          result := input_90;
        WHEN "1011011" =>
          result := input_91;
        WHEN "1011100" =>
          result := input_92;
        WHEN "1011101" =>
          result := input_93;
        WHEN "1011110" =>
          result := input_94;
        WHEN "1011111" =>
          result := input_95;
        WHEN "1100000" =>
          result := input_96;
        WHEN "1100001" =>
          result := input_97;
        WHEN "1100010" =>
          result := input_98;
        WHEN "1100011" =>
          result := input_99;
        WHEN "1100100" =>
          result := input_100;
        WHEN "1100101" =>
          result := input_101;
        WHEN "1100110" =>
          result := input_102;
        WHEN "1100111" =>
          result := input_103;
        WHEN "1101000" =>
          result := input_104;
        WHEN "1101001" =>
          result := input_105;
        WHEN "1101010" =>
          result := input_106;
        WHEN "1101011" =>
          result := input_107;
        WHEN "1101100" =>
          result := input_108;
        WHEN "1101101" =>
          result := input_109;
        WHEN "1101110" =>
          result := input_110;
        WHEN "1101111" =>
          result := input_111;
        WHEN "1110000" =>
          result := input_112;
        WHEN "1110001" =>
          result := input_113;
        WHEN "1110010" =>
          result := input_114;
        WHEN "1110011" =>
          result := input_115;
        WHEN "1110100" =>
          result := input_116;
        WHEN "1110101" =>
          result := input_117;
        WHEN "1110110" =>
          result := input_118;
        WHEN "1110111" =>
          result := input_119;
        WHEN "1111000" =>
          result := input_120;
        WHEN "1111001" =>
          result := input_121;
        WHEN "1111010" =>
          result := input_122;
        WHEN "1111011" =>
          result := input_123;
        WHEN "1111100" =>
          result := input_124;
        WHEN "1111101" =>
          result := input_125;
        WHEN "1111110" =>
          result := input_126;
        WHEN others =>
          result := input_127;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_7_2_2(input_0 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(6 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  input_rsci : work.ccs_in_pkg_v1.ccs_in_v1
    GENERIC MAP(
      rscid => 1,
      width => 4096
      )
    PORT MAP(
      dat => input_rsci_dat,
      idat => input_rsci_idat_1
    );
  input_rsci_dat <= input_rsc_dat;
  input_rsci_idat <= input_rsci_idat_1;

  output_rsci : work.ccs_out_pkg_v1.ccs_out_v1
    GENERIC MAP(
      rscid => 2,
      width => 4096
      )
    PORT MAP(
      idat => output_rsci_idat,
      dat => output_rsci_dat
    );
  output_rsci_idat <= output_rsci_idat_4095_4064 & output_rsci_idat_4063_4032 & output_rsci_idat_4031_4000
      & output_rsci_idat_3999_3968 & output_rsci_idat_3967_3936 & output_rsci_idat_3935_3904
      & output_rsci_idat_3903_3872 & output_rsci_idat_3871_3840 & output_rsci_idat_3839_3808
      & output_rsci_idat_3807_3776 & output_rsci_idat_3775_3744 & output_rsci_idat_3743_3712
      & output_rsci_idat_3711_3680 & output_rsci_idat_3679_3648 & output_rsci_idat_3647_3616
      & output_rsci_idat_3615_3584 & output_rsci_idat_3583_3552 & output_rsci_idat_3551_3520
      & output_rsci_idat_3519_3488 & output_rsci_idat_3487_3456 & output_rsci_idat_3455_3424
      & output_rsci_idat_3423_3392 & output_rsci_idat_3391_3360 & output_rsci_idat_3359_3328
      & output_rsci_idat_3327_3296 & output_rsci_idat_3295_3264 & output_rsci_idat_3263_3232
      & output_rsci_idat_3231_3200 & output_rsci_idat_3199_3168 & output_rsci_idat_3167_3136
      & output_rsci_idat_3135_3104 & output_rsci_idat_3103_3072 & output_rsci_idat_3071_3040
      & output_rsci_idat_3039_3008 & output_rsci_idat_3007_2976 & output_rsci_idat_2975_2944
      & output_rsci_idat_2943_2912 & output_rsci_idat_2911_2880 & output_rsci_idat_2879_2848
      & output_rsci_idat_2847_2816 & output_rsci_idat_2815_2784 & output_rsci_idat_2783_2752
      & output_rsci_idat_2751_2720 & output_rsci_idat_2719_2688 & output_rsci_idat_2687_2656
      & output_rsci_idat_2655_2624 & output_rsci_idat_2623_2592 & output_rsci_idat_2591_2560
      & output_rsci_idat_2559_2528 & output_rsci_idat_2527_2496 & output_rsci_idat_2495_2464
      & output_rsci_idat_2463_2432 & output_rsci_idat_2431_2400 & output_rsci_idat_2399_2368
      & output_rsci_idat_2367_2336 & output_rsci_idat_2335_2304 & output_rsci_idat_2303_2272
      & output_rsci_idat_2271_2240 & output_rsci_idat_2239_2208 & output_rsci_idat_2207_2176
      & output_rsci_idat_2175_2144 & output_rsci_idat_2143_2112 & output_rsci_idat_2111_2080
      & output_rsci_idat_2079_2048 & output_rsci_idat_2047_2016 & output_rsci_idat_2015_1984
      & output_rsci_idat_1983_1952 & output_rsci_idat_1951_1920 & output_rsci_idat_1919_1888
      & output_rsci_idat_1887_1856 & output_rsci_idat_1855_1824 & output_rsci_idat_1823_1792
      & output_rsci_idat_1791_1760 & output_rsci_idat_1759_1728 & output_rsci_idat_1727_1696
      & output_rsci_idat_1695_1664 & output_rsci_idat_1663_1632 & output_rsci_idat_1631_1600
      & output_rsci_idat_1599_1568 & output_rsci_idat_1567_1536 & output_rsci_idat_1535_1504
      & output_rsci_idat_1503_1472 & output_rsci_idat_1471_1440 & output_rsci_idat_1439_1408
      & output_rsci_idat_1407_1376 & output_rsci_idat_1375_1344 & output_rsci_idat_1343_1312
      & output_rsci_idat_1311_1280 & output_rsci_idat_1279_1248 & output_rsci_idat_1247_1216
      & output_rsci_idat_1215_1184 & output_rsci_idat_1183_1152 & output_rsci_idat_1151_1120
      & output_rsci_idat_1119_1088 & output_rsci_idat_1087_1056 & output_rsci_idat_1055_1024
      & output_rsci_idat_1023_992 & output_rsci_idat_991_960 & output_rsci_idat_959_928
      & output_rsci_idat_927_896 & output_rsci_idat_895_864 & output_rsci_idat_863_832
      & output_rsci_idat_831_800 & output_rsci_idat_799_768 & output_rsci_idat_767_736
      & output_rsci_idat_735_704 & output_rsci_idat_703_672 & output_rsci_idat_671_640
      & output_rsci_idat_639_608 & output_rsci_idat_607_576 & output_rsci_idat_575_544
      & output_rsci_idat_543_512 & output_rsci_idat_511_480 & output_rsci_idat_479_448
      & output_rsci_idat_447_416 & output_rsci_idat_415_384 & output_rsci_idat_383_352
      & output_rsci_idat_351_320 & output_rsci_idat_319_288 & output_rsci_idat_287_256
      & output_rsci_idat_255_224 & output_rsci_idat_223_192 & output_rsci_idat_191_160
      & output_rsci_idat_159_128 & output_rsci_idat_127_96 & output_rsci_idat_95_64
      & output_rsci_idat_63_32 & output_rsci_idat_31_0;
  output_rsc_dat <= output_rsci_dat;

  input_rsc_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_output_rsc_triosy_obj_ld_cse,
      lz => input_rsc_triosy_lz
    );
  output_rsc_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_output_rsc_triosy_obj_ld_cse,
      lz => output_rsc_triosy_lz
    );
  fir_core_core_fsm_inst : fir_core_core_fsm
    PORT MAP(
      clk => clk,
      rst => rst,
      fsm_output => fir_core_core_fsm_inst_fsm_output,
      for_C_2_tr0 => fir_core_core_fsm_inst_for_C_2_tr0
    );
  fsm_output <= fir_core_core_fsm_inst_fsm_output;
  fir_core_core_fsm_inst_for_C_2_tr0 <= i_7_0_sva_1(7);

  reg_output_rsc_1_31_output_or_cse <= (fsm_output(3)) OR (fsm_output(0));
  output_output_mux_cse <= MUX_v_32_2_2(output_rsc_1_31_0_lpi_2, for_for_mul_1_cmx_sva_1,
      or_tmp_259);
  for_for_mul_1_cmx_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED'( SIGNED(for_mux_itm)
      * SIGNED'( "01101")), 32));
  for_or_tmp <= ((i_7_0_sva_6_0(0)) AND for_nor_itm) OR ((i_7_0_sva_6_0(1)) AND for_nor_1_itm)
      OR for_equal_tmp_3 OR ((i_7_0_sva_6_0(2)) AND for_nor_3_itm) OR for_equal_tmp_5
      OR for_equal_tmp_6 OR for_equal_tmp_7 OR ((i_7_0_sva_6_0(3)) AND for_nor_7_itm)
      OR for_equal_tmp_9 OR for_equal_tmp_10 OR for_equal_tmp_11 OR for_equal_tmp_12
      OR for_equal_tmp_13 OR for_equal_tmp_14 OR for_equal_tmp_15 OR ((i_7_0_sva_6_0(4))
      AND for_nor_15_itm) OR for_equal_tmp_17 OR for_equal_tmp_18 OR for_equal_tmp_19
      OR for_equal_tmp_20 OR for_equal_tmp_21 OR for_equal_tmp_22 OR for_equal_tmp_23
      OR for_equal_tmp_24 OR for_equal_tmp_25 OR for_equal_tmp_26 OR for_equal_tmp_27
      OR for_equal_tmp_28 OR for_equal_tmp_29 OR for_equal_tmp_30 OR for_equal_tmp_31
      OR ((i_7_0_sva_6_0(5)) AND for_nor_31_itm) OR for_equal_tmp_33 OR for_equal_tmp_34
      OR for_equal_tmp_35 OR for_equal_tmp_36 OR for_equal_tmp_37 OR for_equal_tmp_38
      OR for_equal_tmp_39 OR for_equal_tmp_40 OR for_equal_tmp_41 OR for_equal_tmp_42
      OR for_equal_tmp_43 OR for_equal_tmp_44 OR for_equal_tmp_45 OR for_equal_tmp_46
      OR for_equal_tmp_47 OR for_equal_tmp_48 OR for_equal_tmp_49 OR for_equal_tmp_50
      OR for_equal_tmp_51 OR for_equal_tmp_52 OR for_equal_tmp_53 OR for_equal_tmp_54
      OR for_equal_tmp_55 OR for_equal_tmp_56 OR for_equal_tmp_57 OR for_equal_tmp_58
      OR for_equal_tmp_59 OR for_equal_tmp_60 OR for_equal_tmp_61 OR for_equal_tmp_62
      OR for_equal_tmp_63 OR ((i_7_0_sva_6_0(6)) AND for_nor_62_itm) OR for_equal_tmp_65
      OR for_equal_tmp_66 OR for_equal_tmp_67 OR for_equal_tmp_68 OR for_equal_tmp_69
      OR for_equal_tmp_70 OR for_equal_tmp_71 OR for_equal_tmp_72 OR for_equal_tmp_73
      OR for_equal_tmp_74 OR for_equal_tmp_75 OR for_equal_tmp_76 OR for_equal_tmp_77
      OR for_equal_tmp_78 OR for_equal_tmp_79 OR for_equal_tmp_80 OR for_equal_tmp_81
      OR for_equal_tmp_82 OR for_equal_tmp_83 OR for_equal_tmp_84 OR for_equal_tmp_85
      OR for_equal_tmp_86 OR for_equal_tmp_87 OR for_equal_tmp_88 OR for_equal_tmp_89
      OR for_equal_tmp_90 OR for_equal_tmp_91 OR for_equal_tmp_92 OR for_equal_tmp_93
      OR for_equal_tmp_94 OR for_equal_tmp_95 OR for_equal_tmp_96 OR for_equal_tmp_97
      OR for_equal_tmp_98 OR for_equal_tmp_99 OR for_equal_tmp_100 OR for_equal_tmp_101
      OR for_equal_tmp_102 OR for_equal_tmp_103 OR for_equal_tmp_104 OR for_equal_tmp_105
      OR for_equal_tmp_106 OR for_equal_tmp_107 OR for_equal_tmp_108 OR for_equal_tmp_109
      OR for_equal_tmp_110 OR for_equal_tmp_111 OR for_equal_tmp_112 OR for_equal_tmp_113
      OR for_equal_tmp_114 OR for_equal_tmp_115 OR for_equal_tmp_116 OR for_equal_tmp_117
      OR for_equal_tmp_118 OR for_equal_tmp_119 OR for_equal_tmp_120 OR for_equal_tmp_121
      OR for_equal_tmp_122 OR for_equal_tmp_123 OR for_equal_tmp_124 OR for_equal_tmp_125
      OR for_equal_tmp_126 OR for_equal_tmp_127;
  or_dcpl_330 <= NOT((i_7_0_sva_6_0(0)) AND for_nor_itm);
  or_dcpl_331 <= NOT((i_7_0_sva_6_0(1)) AND for_nor_1_itm);
  or_dcpl_332 <= NOT((i_7_0_sva_6_0(2)) AND for_nor_3_itm);
  or_dcpl_333 <= NOT((i_7_0_sva_6_0(3)) AND for_nor_7_itm);
  or_dcpl_334 <= NOT((i_7_0_sva_6_0(4)) AND for_nor_15_itm);
  or_dcpl_335 <= NOT((i_7_0_sva_6_0(5)) AND for_nor_31_itm);
  or_dcpl_336 <= NOT(for_nor_62_itm AND (i_7_0_sva_6_0(6)));
  or_tmp_259 <= (NOT for_or_tmp) AND (fsm_output(2));
  or_tmp_643 <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00"));
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsc_1_31_0_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_63_32_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_95_64_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_127_96_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_159_128_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_191_160_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_223_192_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_255_224_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_287_256_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_319_288_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_351_320_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_383_352_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_415_384_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_447_416_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_479_448_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_511_480_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_543_512_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_575_544_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_607_576_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_639_608_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_671_640_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_703_672_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_735_704_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_767_736_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_799_768_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_831_800_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_863_832_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_895_864_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_927_896_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_959_928_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_991_960_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_1023_992_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_1055_1024_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_1087_1056_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_1119_1088_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_1151_1120_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_1183_1152_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_1215_1184_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_1247_1216_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_1279_1248_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_1311_1280_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_1343_1312_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_1375_1344_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_1407_1376_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_1439_1408_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_1471_1440_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_1503_1472_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_1535_1504_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_1567_1536_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_1599_1568_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_1631_1600_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_1663_1632_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_1695_1664_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_1727_1696_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_1759_1728_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_1791_1760_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_1823_1792_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_1855_1824_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_1887_1856_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_1919_1888_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_1951_1920_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_1983_1952_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_2015_1984_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_2047_2016_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_2079_2048_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_2111_2080_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_2143_2112_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_2175_2144_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_2207_2176_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_2239_2208_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_2271_2240_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_2303_2272_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_2335_2304_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_2367_2336_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_2399_2368_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_2431_2400_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_2463_2432_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_2495_2464_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_2527_2496_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_2559_2528_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_2591_2560_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_2623_2592_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_2655_2624_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_2687_2656_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_2719_2688_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_2751_2720_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_2783_2752_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_2815_2784_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_2847_2816_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_2879_2848_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_2911_2880_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_2943_2912_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_2975_2944_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_3007_2976_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_3039_3008_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_3071_3040_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_3103_3072_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_3135_3104_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_3167_3136_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_3199_3168_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_3231_3200_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_3263_3232_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_3295_3264_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_3327_3296_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_3359_3328_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_3391_3360_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_3423_3392_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_3455_3424_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_3487_3456_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_3519_3488_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_3551_3520_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_3583_3552_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_3615_3584_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_3647_3616_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_3679_3648_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_3711_3680_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_3743_3712_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_3775_3744_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_3807_3776_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_3839_3808_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_3871_3840_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_3903_3872_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_3935_3904_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_3967_3936_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_3999_3968_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_4031_4000_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_4063_4032_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        output_rsc_1_4095_4064_lpi_2 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        i_7_0_sva_6_0 <= STD_LOGIC_VECTOR'( "0000000");
      ELSIF ( reg_output_rsc_1_31_output_or_cse = '1' ) THEN
        output_rsc_1_31_0_lpi_2 <= for_io_read_output_rsc_sdt_31_0_lpi_2_dfm;
        output_rsc_1_63_32_lpi_2 <= for_io_read_output_rsc_sdt_63_32_lpi_2_dfm;
        output_rsc_1_95_64_lpi_2 <= for_io_read_output_rsc_sdt_95_64_lpi_2_dfm;
        output_rsc_1_127_96_lpi_2 <= for_io_read_output_rsc_sdt_127_96_lpi_2_dfm;
        output_rsc_1_159_128_lpi_2 <= for_io_read_output_rsc_sdt_159_128_lpi_2_dfm;
        output_rsc_1_191_160_lpi_2 <= for_io_read_output_rsc_sdt_191_160_lpi_2_dfm;
        output_rsc_1_223_192_lpi_2 <= for_io_read_output_rsc_sdt_223_192_lpi_2_dfm;
        output_rsc_1_255_224_lpi_2 <= for_io_read_output_rsc_sdt_255_224_lpi_2_dfm;
        output_rsc_1_287_256_lpi_2 <= for_io_read_output_rsc_sdt_287_256_lpi_2_dfm;
        output_rsc_1_319_288_lpi_2 <= for_io_read_output_rsc_sdt_319_288_lpi_2_dfm;
        output_rsc_1_351_320_lpi_2 <= for_io_read_output_rsc_sdt_351_320_lpi_2_dfm;
        output_rsc_1_383_352_lpi_2 <= for_io_read_output_rsc_sdt_383_352_lpi_2_dfm;
        output_rsc_1_415_384_lpi_2 <= for_io_read_output_rsc_sdt_415_384_lpi_2_dfm;
        output_rsc_1_447_416_lpi_2 <= for_io_read_output_rsc_sdt_447_416_lpi_2_dfm;
        output_rsc_1_479_448_lpi_2 <= for_io_read_output_rsc_sdt_479_448_lpi_2_dfm;
        output_rsc_1_511_480_lpi_2 <= for_io_read_output_rsc_sdt_511_480_lpi_2_dfm;
        output_rsc_1_543_512_lpi_2 <= for_io_read_output_rsc_sdt_543_512_lpi_2_dfm;
        output_rsc_1_575_544_lpi_2 <= for_io_read_output_rsc_sdt_575_544_lpi_2_dfm;
        output_rsc_1_607_576_lpi_2 <= for_io_read_output_rsc_sdt_607_576_lpi_2_dfm;
        output_rsc_1_639_608_lpi_2 <= for_io_read_output_rsc_sdt_639_608_lpi_2_dfm;
        output_rsc_1_671_640_lpi_2 <= for_io_read_output_rsc_sdt_671_640_lpi_2_dfm;
        output_rsc_1_703_672_lpi_2 <= for_io_read_output_rsc_sdt_703_672_lpi_2_dfm;
        output_rsc_1_735_704_lpi_2 <= for_io_read_output_rsc_sdt_735_704_lpi_2_dfm;
        output_rsc_1_767_736_lpi_2 <= for_io_read_output_rsc_sdt_767_736_lpi_2_dfm;
        output_rsc_1_799_768_lpi_2 <= for_io_read_output_rsc_sdt_799_768_lpi_2_dfm;
        output_rsc_1_831_800_lpi_2 <= for_io_read_output_rsc_sdt_831_800_lpi_2_dfm;
        output_rsc_1_863_832_lpi_2 <= for_io_read_output_rsc_sdt_863_832_lpi_2_dfm;
        output_rsc_1_895_864_lpi_2 <= for_io_read_output_rsc_sdt_895_864_lpi_2_dfm;
        output_rsc_1_927_896_lpi_2 <= for_io_read_output_rsc_sdt_927_896_lpi_2_dfm;
        output_rsc_1_959_928_lpi_2 <= for_io_read_output_rsc_sdt_959_928_lpi_2_dfm;
        output_rsc_1_991_960_lpi_2 <= for_io_read_output_rsc_sdt_991_960_lpi_2_dfm;
        output_rsc_1_1023_992_lpi_2 <= for_io_read_output_rsc_sdt_1023_992_lpi_2_dfm;
        output_rsc_1_1055_1024_lpi_2 <= for_io_read_output_rsc_sdt_1055_1024_lpi_2_dfm;
        output_rsc_1_1087_1056_lpi_2 <= for_io_read_output_rsc_sdt_1087_1056_lpi_2_dfm;
        output_rsc_1_1119_1088_lpi_2 <= for_io_read_output_rsc_sdt_1119_1088_lpi_2_dfm;
        output_rsc_1_1151_1120_lpi_2 <= for_io_read_output_rsc_sdt_1151_1120_lpi_2_dfm;
        output_rsc_1_1183_1152_lpi_2 <= for_io_read_output_rsc_sdt_1183_1152_lpi_2_dfm;
        output_rsc_1_1215_1184_lpi_2 <= for_io_read_output_rsc_sdt_1215_1184_lpi_2_dfm;
        output_rsc_1_1247_1216_lpi_2 <= for_io_read_output_rsc_sdt_1247_1216_lpi_2_dfm;
        output_rsc_1_1279_1248_lpi_2 <= for_io_read_output_rsc_sdt_1279_1248_lpi_2_dfm;
        output_rsc_1_1311_1280_lpi_2 <= for_io_read_output_rsc_sdt_1311_1280_lpi_2_dfm;
        output_rsc_1_1343_1312_lpi_2 <= for_io_read_output_rsc_sdt_1343_1312_lpi_2_dfm;
        output_rsc_1_1375_1344_lpi_2 <= for_io_read_output_rsc_sdt_1375_1344_lpi_2_dfm;
        output_rsc_1_1407_1376_lpi_2 <= for_io_read_output_rsc_sdt_1407_1376_lpi_2_dfm;
        output_rsc_1_1439_1408_lpi_2 <= for_io_read_output_rsc_sdt_1439_1408_lpi_2_dfm;
        output_rsc_1_1471_1440_lpi_2 <= for_io_read_output_rsc_sdt_1471_1440_lpi_2_dfm;
        output_rsc_1_1503_1472_lpi_2 <= for_io_read_output_rsc_sdt_1503_1472_lpi_2_dfm;
        output_rsc_1_1535_1504_lpi_2 <= for_io_read_output_rsc_sdt_1535_1504_lpi_2_dfm;
        output_rsc_1_1567_1536_lpi_2 <= for_io_read_output_rsc_sdt_1567_1536_lpi_2_dfm;
        output_rsc_1_1599_1568_lpi_2 <= for_io_read_output_rsc_sdt_1599_1568_lpi_2_dfm;
        output_rsc_1_1631_1600_lpi_2 <= for_io_read_output_rsc_sdt_1631_1600_lpi_2_dfm;
        output_rsc_1_1663_1632_lpi_2 <= for_io_read_output_rsc_sdt_1663_1632_lpi_2_dfm;
        output_rsc_1_1695_1664_lpi_2 <= for_io_read_output_rsc_sdt_1695_1664_lpi_2_dfm;
        output_rsc_1_1727_1696_lpi_2 <= for_io_read_output_rsc_sdt_1727_1696_lpi_2_dfm;
        output_rsc_1_1759_1728_lpi_2 <= for_io_read_output_rsc_sdt_1759_1728_lpi_2_dfm;
        output_rsc_1_1791_1760_lpi_2 <= for_io_read_output_rsc_sdt_1791_1760_lpi_2_dfm;
        output_rsc_1_1823_1792_lpi_2 <= for_io_read_output_rsc_sdt_1823_1792_lpi_2_dfm;
        output_rsc_1_1855_1824_lpi_2 <= for_io_read_output_rsc_sdt_1855_1824_lpi_2_dfm;
        output_rsc_1_1887_1856_lpi_2 <= for_io_read_output_rsc_sdt_1887_1856_lpi_2_dfm;
        output_rsc_1_1919_1888_lpi_2 <= for_io_read_output_rsc_sdt_1919_1888_lpi_2_dfm;
        output_rsc_1_1951_1920_lpi_2 <= for_io_read_output_rsc_sdt_1951_1920_lpi_2_dfm;
        output_rsc_1_1983_1952_lpi_2 <= for_io_read_output_rsc_sdt_1983_1952_lpi_2_dfm;
        output_rsc_1_2015_1984_lpi_2 <= for_io_read_output_rsc_sdt_2015_1984_lpi_2_dfm;
        output_rsc_1_2047_2016_lpi_2 <= for_io_read_output_rsc_sdt_2047_2016_lpi_2_dfm;
        output_rsc_1_2079_2048_lpi_2 <= for_io_read_output_rsc_sdt_2079_2048_lpi_2_dfm;
        output_rsc_1_2111_2080_lpi_2 <= for_io_read_output_rsc_sdt_2111_2080_lpi_2_dfm;
        output_rsc_1_2143_2112_lpi_2 <= for_io_read_output_rsc_sdt_2143_2112_lpi_2_dfm;
        output_rsc_1_2175_2144_lpi_2 <= for_io_read_output_rsc_sdt_2175_2144_lpi_2_dfm;
        output_rsc_1_2207_2176_lpi_2 <= for_io_read_output_rsc_sdt_2207_2176_lpi_2_dfm;
        output_rsc_1_2239_2208_lpi_2 <= for_io_read_output_rsc_sdt_2239_2208_lpi_2_dfm;
        output_rsc_1_2271_2240_lpi_2 <= for_io_read_output_rsc_sdt_2271_2240_lpi_2_dfm;
        output_rsc_1_2303_2272_lpi_2 <= for_io_read_output_rsc_sdt_2303_2272_lpi_2_dfm;
        output_rsc_1_2335_2304_lpi_2 <= for_io_read_output_rsc_sdt_2335_2304_lpi_2_dfm;
        output_rsc_1_2367_2336_lpi_2 <= for_io_read_output_rsc_sdt_2367_2336_lpi_2_dfm;
        output_rsc_1_2399_2368_lpi_2 <= for_io_read_output_rsc_sdt_2399_2368_lpi_2_dfm;
        output_rsc_1_2431_2400_lpi_2 <= for_io_read_output_rsc_sdt_2431_2400_lpi_2_dfm;
        output_rsc_1_2463_2432_lpi_2 <= for_io_read_output_rsc_sdt_2463_2432_lpi_2_dfm;
        output_rsc_1_2495_2464_lpi_2 <= for_io_read_output_rsc_sdt_2495_2464_lpi_2_dfm;
        output_rsc_1_2527_2496_lpi_2 <= for_io_read_output_rsc_sdt_2527_2496_lpi_2_dfm;
        output_rsc_1_2559_2528_lpi_2 <= for_io_read_output_rsc_sdt_2559_2528_lpi_2_dfm;
        output_rsc_1_2591_2560_lpi_2 <= for_io_read_output_rsc_sdt_2591_2560_lpi_2_dfm;
        output_rsc_1_2623_2592_lpi_2 <= for_io_read_output_rsc_sdt_2623_2592_lpi_2_dfm;
        output_rsc_1_2655_2624_lpi_2 <= for_io_read_output_rsc_sdt_2655_2624_lpi_2_dfm;
        output_rsc_1_2687_2656_lpi_2 <= for_io_read_output_rsc_sdt_2687_2656_lpi_2_dfm;
        output_rsc_1_2719_2688_lpi_2 <= for_io_read_output_rsc_sdt_2719_2688_lpi_2_dfm;
        output_rsc_1_2751_2720_lpi_2 <= for_io_read_output_rsc_sdt_2751_2720_lpi_2_dfm;
        output_rsc_1_2783_2752_lpi_2 <= for_io_read_output_rsc_sdt_2783_2752_lpi_2_dfm;
        output_rsc_1_2815_2784_lpi_2 <= for_io_read_output_rsc_sdt_2815_2784_lpi_2_dfm;
        output_rsc_1_2847_2816_lpi_2 <= for_io_read_output_rsc_sdt_2847_2816_lpi_2_dfm;
        output_rsc_1_2879_2848_lpi_2 <= for_io_read_output_rsc_sdt_2879_2848_lpi_2_dfm;
        output_rsc_1_2911_2880_lpi_2 <= for_io_read_output_rsc_sdt_2911_2880_lpi_2_dfm;
        output_rsc_1_2943_2912_lpi_2 <= for_io_read_output_rsc_sdt_2943_2912_lpi_2_dfm;
        output_rsc_1_2975_2944_lpi_2 <= for_io_read_output_rsc_sdt_2975_2944_lpi_2_dfm;
        output_rsc_1_3007_2976_lpi_2 <= for_io_read_output_rsc_sdt_3007_2976_lpi_2_dfm;
        output_rsc_1_3039_3008_lpi_2 <= for_io_read_output_rsc_sdt_3039_3008_lpi_2_dfm;
        output_rsc_1_3071_3040_lpi_2 <= for_io_read_output_rsc_sdt_3071_3040_lpi_2_dfm;
        output_rsc_1_3103_3072_lpi_2 <= for_io_read_output_rsc_sdt_3103_3072_lpi_2_dfm;
        output_rsc_1_3135_3104_lpi_2 <= for_io_read_output_rsc_sdt_3135_3104_lpi_2_dfm;
        output_rsc_1_3167_3136_lpi_2 <= for_io_read_output_rsc_sdt_3167_3136_lpi_2_dfm;
        output_rsc_1_3199_3168_lpi_2 <= for_io_read_output_rsc_sdt_3199_3168_lpi_2_dfm;
        output_rsc_1_3231_3200_lpi_2 <= for_io_read_output_rsc_sdt_3231_3200_lpi_2_dfm;
        output_rsc_1_3263_3232_lpi_2 <= for_io_read_output_rsc_sdt_3263_3232_lpi_2_dfm;
        output_rsc_1_3295_3264_lpi_2 <= for_io_read_output_rsc_sdt_3295_3264_lpi_2_dfm;
        output_rsc_1_3327_3296_lpi_2 <= for_io_read_output_rsc_sdt_3327_3296_lpi_2_dfm;
        output_rsc_1_3359_3328_lpi_2 <= for_io_read_output_rsc_sdt_3359_3328_lpi_2_dfm;
        output_rsc_1_3391_3360_lpi_2 <= for_io_read_output_rsc_sdt_3391_3360_lpi_2_dfm;
        output_rsc_1_3423_3392_lpi_2 <= for_io_read_output_rsc_sdt_3423_3392_lpi_2_dfm;
        output_rsc_1_3455_3424_lpi_2 <= for_io_read_output_rsc_sdt_3455_3424_lpi_2_dfm;
        output_rsc_1_3487_3456_lpi_2 <= for_io_read_output_rsc_sdt_3487_3456_lpi_2_dfm;
        output_rsc_1_3519_3488_lpi_2 <= for_io_read_output_rsc_sdt_3519_3488_lpi_2_dfm;
        output_rsc_1_3551_3520_lpi_2 <= for_io_read_output_rsc_sdt_3551_3520_lpi_2_dfm;
        output_rsc_1_3583_3552_lpi_2 <= for_io_read_output_rsc_sdt_3583_3552_lpi_2_dfm;
        output_rsc_1_3615_3584_lpi_2 <= for_io_read_output_rsc_sdt_3615_3584_lpi_2_dfm;
        output_rsc_1_3647_3616_lpi_2 <= for_io_read_output_rsc_sdt_3647_3616_lpi_2_dfm;
        output_rsc_1_3679_3648_lpi_2 <= for_io_read_output_rsc_sdt_3679_3648_lpi_2_dfm;
        output_rsc_1_3711_3680_lpi_2 <= for_io_read_output_rsc_sdt_3711_3680_lpi_2_dfm;
        output_rsc_1_3743_3712_lpi_2 <= for_io_read_output_rsc_sdt_3743_3712_lpi_2_dfm;
        output_rsc_1_3775_3744_lpi_2 <= for_io_read_output_rsc_sdt_3775_3744_lpi_2_dfm;
        output_rsc_1_3807_3776_lpi_2 <= for_io_read_output_rsc_sdt_3807_3776_lpi_2_dfm;
        output_rsc_1_3839_3808_lpi_2 <= for_io_read_output_rsc_sdt_3839_3808_lpi_2_dfm;
        output_rsc_1_3871_3840_lpi_2 <= for_io_read_output_rsc_sdt_3871_3840_lpi_2_dfm;
        output_rsc_1_3903_3872_lpi_2 <= for_io_read_output_rsc_sdt_3903_3872_lpi_2_dfm;
        output_rsc_1_3935_3904_lpi_2 <= for_io_read_output_rsc_sdt_3935_3904_lpi_2_dfm;
        output_rsc_1_3967_3936_lpi_2 <= for_io_read_output_rsc_sdt_3967_3936_lpi_2_dfm;
        output_rsc_1_3999_3968_lpi_2 <= for_io_read_output_rsc_sdt_3999_3968_lpi_2_dfm;
        output_rsc_1_4031_4000_lpi_2 <= for_io_read_output_rsc_sdt_4031_4000_lpi_2_dfm;
        output_rsc_1_4063_4032_lpi_2 <= for_io_read_output_rsc_sdt_4063_4032_lpi_2_dfm;
        output_rsc_1_4095_4064_lpi_2 <= for_io_read_output_rsc_sdt_4095_4064_lpi_2_dfm;
        i_7_0_sva_6_0 <= MUX_v_7_2_2(STD_LOGIC_VECTOR'("0000000"), (i_7_0_sva_1(6
            DOWNTO 0)), (fsm_output(3)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_31_0 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( ((for_or_tmp AND (fsm_output(2))) OR or_tmp_259) = '1' ) THEN
        output_rsci_idat_31_0 <= output_output_mux_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_63_32 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_63_32 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_63_32_lpi_2,
            and_660_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_95_64 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_95_64 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_95_64_lpi_2,
            and_666_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_127_96 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_127_96 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_127_96_lpi_2,
            and_672_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_159_128 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_159_128 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_159_128_lpi_2,
            and_678_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_191_160 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_191_160 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_191_160_lpi_2,
            and_684_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_223_192 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_223_192 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_223_192_lpi_2,
            and_690_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_255_224 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_255_224 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_255_224_lpi_2,
            and_696_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_287_256 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_287_256 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_287_256_lpi_2,
            and_702_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_319_288 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_319_288 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_319_288_lpi_2,
            and_708_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_351_320 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_351_320 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_351_320_lpi_2,
            and_714_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_383_352 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_383_352 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_383_352_lpi_2,
            and_720_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_415_384 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_415_384 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_415_384_lpi_2,
            and_726_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_447_416 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_447_416 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_447_416_lpi_2,
            and_732_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_479_448 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_479_448 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_479_448_lpi_2,
            and_738_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_511_480 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_511_480 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_511_480_lpi_2,
            and_744_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_543_512 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_543_512 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_543_512_lpi_2,
            and_750_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_575_544 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_575_544 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_575_544_lpi_2,
            and_756_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_607_576 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_607_576 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_607_576_lpi_2,
            and_762_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_639_608 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_639_608 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_639_608_lpi_2,
            and_768_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_671_640 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_671_640 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_671_640_lpi_2,
            and_774_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_703_672 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_703_672 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_703_672_lpi_2,
            and_780_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_735_704 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_735_704 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_735_704_lpi_2,
            and_786_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_767_736 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_767_736 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_767_736_lpi_2,
            and_792_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_799_768 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_799_768 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_799_768_lpi_2,
            and_798_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_831_800 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_831_800 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_831_800_lpi_2,
            and_804_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_863_832 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_863_832 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_863_832_lpi_2,
            and_810_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_895_864 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_895_864 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_895_864_lpi_2,
            and_816_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_927_896 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_927_896 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_927_896_lpi_2,
            and_822_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_959_928 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_959_928 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_959_928_lpi_2,
            and_828_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_991_960 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_991_960 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_991_960_lpi_2,
            and_834_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_1023_992 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_1023_992 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1023_992_lpi_2,
            and_840_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_1055_1024 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_1055_1024 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1055_1024_lpi_2,
            and_846_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_1087_1056 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_1087_1056 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1087_1056_lpi_2,
            and_852_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_1119_1088 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_1119_1088 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1119_1088_lpi_2,
            and_858_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_1151_1120 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_1151_1120 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1151_1120_lpi_2,
            and_864_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_1183_1152 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_1183_1152 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1183_1152_lpi_2,
            and_870_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_1215_1184 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_1215_1184 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1215_1184_lpi_2,
            and_876_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_1247_1216 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_1247_1216 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1247_1216_lpi_2,
            and_882_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_1279_1248 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_1279_1248 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1279_1248_lpi_2,
            and_888_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_1311_1280 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_1311_1280 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1311_1280_lpi_2,
            and_894_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_1343_1312 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_1343_1312 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1343_1312_lpi_2,
            and_900_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_1375_1344 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_1375_1344 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1375_1344_lpi_2,
            and_906_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_1407_1376 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_1407_1376 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1407_1376_lpi_2,
            and_912_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_1439_1408 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_1439_1408 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1439_1408_lpi_2,
            and_918_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_1471_1440 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_1471_1440 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1471_1440_lpi_2,
            and_924_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_1503_1472 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_1503_1472 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1503_1472_lpi_2,
            and_930_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_1535_1504 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_1535_1504 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1535_1504_lpi_2,
            and_936_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_1567_1536 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_1567_1536 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1567_1536_lpi_2,
            and_942_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_1599_1568 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_1599_1568 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1599_1568_lpi_2,
            and_948_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_1631_1600 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_1631_1600 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1631_1600_lpi_2,
            and_954_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_1663_1632 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_1663_1632 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1663_1632_lpi_2,
            and_960_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_1695_1664 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_1695_1664 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1695_1664_lpi_2,
            and_966_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_1727_1696 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_1727_1696 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1727_1696_lpi_2,
            and_972_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_1759_1728 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_1759_1728 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1759_1728_lpi_2,
            and_978_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_1791_1760 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_1791_1760 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1791_1760_lpi_2,
            and_984_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_1823_1792 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_1823_1792 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1823_1792_lpi_2,
            and_990_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_1855_1824 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_1855_1824 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1855_1824_lpi_2,
            and_996_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_1887_1856 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_1887_1856 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1887_1856_lpi_2,
            and_1002_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_1919_1888 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_1919_1888 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1919_1888_lpi_2,
            and_1008_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_1951_1920 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_1951_1920 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1951_1920_lpi_2,
            and_1014_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_1983_1952 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_1983_1952 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1983_1952_lpi_2,
            and_1020_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_2015_1984 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_2015_1984 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2015_1984_lpi_2,
            and_1026_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_2047_2016 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_2047_2016 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2047_2016_lpi_2,
            and_1032_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_2079_2048 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_2079_2048 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2079_2048_lpi_2,
            and_1038_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_2111_2080 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_2111_2080 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2111_2080_lpi_2,
            and_1044_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_2143_2112 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_2143_2112 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2143_2112_lpi_2,
            and_1050_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_2175_2144 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_2175_2144 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2175_2144_lpi_2,
            and_1056_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_2207_2176 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_2207_2176 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2207_2176_lpi_2,
            and_1062_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_2239_2208 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_2239_2208 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2239_2208_lpi_2,
            and_1068_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_2271_2240 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_2271_2240 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2271_2240_lpi_2,
            and_1074_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_2303_2272 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_2303_2272 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2303_2272_lpi_2,
            and_1080_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_2335_2304 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_2335_2304 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2335_2304_lpi_2,
            and_1086_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_2367_2336 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_2367_2336 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2367_2336_lpi_2,
            and_1092_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_2399_2368 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_2399_2368 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2399_2368_lpi_2,
            and_1098_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_2431_2400 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_2431_2400 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2431_2400_lpi_2,
            and_1104_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_2463_2432 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_2463_2432 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2463_2432_lpi_2,
            and_1110_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_2495_2464 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_2495_2464 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2495_2464_lpi_2,
            and_1116_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_2527_2496 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_2527_2496 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2527_2496_lpi_2,
            and_1122_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_2559_2528 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_2559_2528 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2559_2528_lpi_2,
            and_1128_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_2591_2560 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_2591_2560 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2591_2560_lpi_2,
            and_1134_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_2623_2592 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_2623_2592 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2623_2592_lpi_2,
            and_1140_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_2655_2624 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_2655_2624 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2655_2624_lpi_2,
            and_1146_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_2687_2656 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_2687_2656 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2687_2656_lpi_2,
            and_1152_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_2719_2688 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_2719_2688 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2719_2688_lpi_2,
            and_1158_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_2751_2720 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_2751_2720 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2751_2720_lpi_2,
            and_1164_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_2783_2752 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_2783_2752 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2783_2752_lpi_2,
            and_1170_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_2815_2784 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_2815_2784 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2815_2784_lpi_2,
            and_1176_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_2847_2816 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_2847_2816 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2847_2816_lpi_2,
            and_1182_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_2879_2848 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_2879_2848 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2879_2848_lpi_2,
            and_1188_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_2911_2880 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_2911_2880 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2911_2880_lpi_2,
            and_1194_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_2943_2912 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_2943_2912 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2943_2912_lpi_2,
            and_1200_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_2975_2944 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_2975_2944 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2975_2944_lpi_2,
            and_1206_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_3007_2976 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_3007_2976 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3007_2976_lpi_2,
            and_1212_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_3039_3008 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_3039_3008 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3039_3008_lpi_2,
            and_1218_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_3071_3040 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_3071_3040 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3071_3040_lpi_2,
            and_1224_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_3103_3072 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_3103_3072 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3103_3072_lpi_2,
            and_1230_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_3135_3104 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_3135_3104 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3135_3104_lpi_2,
            and_1236_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_3167_3136 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_3167_3136 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3167_3136_lpi_2,
            and_1242_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_3199_3168 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_3199_3168 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3199_3168_lpi_2,
            and_1248_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_3231_3200 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_3231_3200 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3231_3200_lpi_2,
            and_1254_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_3263_3232 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_3263_3232 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3263_3232_lpi_2,
            and_1260_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_3295_3264 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_3295_3264 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3295_3264_lpi_2,
            and_1266_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_3327_3296 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_3327_3296 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3327_3296_lpi_2,
            and_1272_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_3359_3328 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_3359_3328 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3359_3328_lpi_2,
            and_1278_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_3391_3360 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_3391_3360 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3391_3360_lpi_2,
            and_1284_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_3423_3392 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_3423_3392 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3423_3392_lpi_2,
            and_1290_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_3455_3424 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_3455_3424 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3455_3424_lpi_2,
            and_1296_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_3487_3456 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_3487_3456 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3487_3456_lpi_2,
            and_1302_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_3519_3488 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_3519_3488 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3519_3488_lpi_2,
            and_1308_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_3551_3520 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_3551_3520 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3551_3520_lpi_2,
            and_1314_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_3583_3552 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_3583_3552 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3583_3552_lpi_2,
            and_1320_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_3615_3584 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_3615_3584 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3615_3584_lpi_2,
            and_1326_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_3647_3616 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_3647_3616 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3647_3616_lpi_2,
            and_1332_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_3679_3648 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_3679_3648 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3679_3648_lpi_2,
            and_1338_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_3711_3680 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_3711_3680 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3711_3680_lpi_2,
            and_1344_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_3743_3712 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_3743_3712 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3743_3712_lpi_2,
            and_1350_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_3775_3744 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_3775_3744 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3775_3744_lpi_2,
            and_1356_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_3807_3776 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_3807_3776 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3807_3776_lpi_2,
            and_1362_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_3839_3808 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_3839_3808 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3839_3808_lpi_2,
            and_1368_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_3871_3840 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_3871_3840 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3871_3840_lpi_2,
            and_1374_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_3903_3872 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_3903_3872 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3903_3872_lpi_2,
            and_1380_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_3935_3904 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_3935_3904 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3935_3904_lpi_2,
            and_1386_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_3967_3936 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_3967_3936 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3967_3936_lpi_2,
            and_1392_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_3999_3968 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_3999_3968 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3999_3968_lpi_2,
            and_1398_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_4031_4000 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_4031_4000 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_4031_4000_lpi_2,
            and_1404_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_4063_4032 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_4063_4032 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_4063_4032_lpi_2,
            and_1410_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat_4095_4064 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( (fsm_output(2)) = '1' ) THEN
        output_rsci_idat_4095_4064 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_4095_4064_lpi_2,
            and_1416_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_output_rsc_triosy_obj_ld_cse <= '0';
        for_equal_tmp_3 <= '0';
        for_equal_tmp_5 <= '0';
        for_equal_tmp_6 <= '0';
        for_equal_tmp_7 <= '0';
        for_equal_tmp_9 <= '0';
        for_equal_tmp_10 <= '0';
        for_equal_tmp_11 <= '0';
        for_equal_tmp_12 <= '0';
        for_equal_tmp_13 <= '0';
        for_equal_tmp_14 <= '0';
        for_equal_tmp_15 <= '0';
        for_equal_tmp_17 <= '0';
        for_equal_tmp_18 <= '0';
        for_equal_tmp_19 <= '0';
        for_equal_tmp_20 <= '0';
        for_equal_tmp_21 <= '0';
        for_equal_tmp_22 <= '0';
        for_equal_tmp_23 <= '0';
        for_equal_tmp_24 <= '0';
        for_equal_tmp_25 <= '0';
        for_equal_tmp_26 <= '0';
        for_equal_tmp_27 <= '0';
        for_equal_tmp_28 <= '0';
        for_equal_tmp_29 <= '0';
        for_equal_tmp_30 <= '0';
        for_equal_tmp_31 <= '0';
        for_equal_tmp_33 <= '0';
        for_equal_tmp_34 <= '0';
        for_equal_tmp_35 <= '0';
        for_equal_tmp_36 <= '0';
        for_equal_tmp_37 <= '0';
        for_equal_tmp_38 <= '0';
        for_equal_tmp_39 <= '0';
        for_equal_tmp_40 <= '0';
        for_equal_tmp_41 <= '0';
        for_equal_tmp_42 <= '0';
        for_equal_tmp_43 <= '0';
        for_equal_tmp_44 <= '0';
        for_equal_tmp_45 <= '0';
        for_equal_tmp_46 <= '0';
        for_equal_tmp_47 <= '0';
        for_equal_tmp_48 <= '0';
        for_equal_tmp_49 <= '0';
        for_equal_tmp_50 <= '0';
        for_equal_tmp_51 <= '0';
        for_equal_tmp_52 <= '0';
        for_equal_tmp_53 <= '0';
        for_equal_tmp_54 <= '0';
        for_equal_tmp_55 <= '0';
        for_equal_tmp_56 <= '0';
        for_equal_tmp_57 <= '0';
        for_equal_tmp_58 <= '0';
        for_equal_tmp_59 <= '0';
        for_equal_tmp_60 <= '0';
        for_equal_tmp_61 <= '0';
        for_equal_tmp_62 <= '0';
        for_equal_tmp_63 <= '0';
        for_equal_tmp_65 <= '0';
        for_equal_tmp_66 <= '0';
        for_equal_tmp_67 <= '0';
        for_equal_tmp_68 <= '0';
        for_equal_tmp_69 <= '0';
        for_equal_tmp_70 <= '0';
        for_equal_tmp_71 <= '0';
        for_equal_tmp_72 <= '0';
        for_equal_tmp_73 <= '0';
        for_equal_tmp_74 <= '0';
        for_equal_tmp_75 <= '0';
        for_equal_tmp_76 <= '0';
        for_equal_tmp_77 <= '0';
        for_equal_tmp_78 <= '0';
        for_equal_tmp_79 <= '0';
        for_equal_tmp_80 <= '0';
        for_equal_tmp_81 <= '0';
        for_equal_tmp_82 <= '0';
        for_equal_tmp_83 <= '0';
        for_equal_tmp_84 <= '0';
        for_equal_tmp_85 <= '0';
        for_equal_tmp_86 <= '0';
        for_equal_tmp_87 <= '0';
        for_equal_tmp_88 <= '0';
        for_equal_tmp_89 <= '0';
        for_equal_tmp_90 <= '0';
        for_equal_tmp_91 <= '0';
        for_equal_tmp_92 <= '0';
        for_equal_tmp_93 <= '0';
        for_equal_tmp_94 <= '0';
        for_equal_tmp_95 <= '0';
        for_equal_tmp_96 <= '0';
        for_equal_tmp_97 <= '0';
        for_equal_tmp_98 <= '0';
        for_equal_tmp_99 <= '0';
        for_equal_tmp_100 <= '0';
        for_equal_tmp_101 <= '0';
        for_equal_tmp_102 <= '0';
        for_equal_tmp_103 <= '0';
        for_equal_tmp_104 <= '0';
        for_equal_tmp_105 <= '0';
        for_equal_tmp_106 <= '0';
        for_equal_tmp_107 <= '0';
        for_equal_tmp_108 <= '0';
        for_equal_tmp_109 <= '0';
        for_equal_tmp_110 <= '0';
        for_equal_tmp_111 <= '0';
        for_equal_tmp_112 <= '0';
        for_equal_tmp_113 <= '0';
        for_equal_tmp_114 <= '0';
        for_equal_tmp_115 <= '0';
        for_equal_tmp_116 <= '0';
        for_equal_tmp_117 <= '0';
        for_equal_tmp_118 <= '0';
        for_equal_tmp_119 <= '0';
        for_equal_tmp_120 <= '0';
        for_equal_tmp_121 <= '0';
        for_equal_tmp_122 <= '0';
        for_equal_tmp_123 <= '0';
        for_equal_tmp_124 <= '0';
        for_equal_tmp_125 <= '0';
        for_equal_tmp_126 <= '0';
        for_equal_tmp_127 <= '0';
        for_nor_62_itm <= '0';
        for_nor_31_itm <= '0';
        for_nor_15_itm <= '0';
        for_nor_7_itm <= '0';
        for_nor_3_itm <= '0';
        for_nor_1_itm <= '0';
        for_nor_itm <= '0';
        for_mux_itm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSE
        reg_output_rsc_triosy_obj_ld_cse <= (i_7_0_sva_1(7)) AND (fsm_output(3));
        for_equal_tmp_3 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0000011"));
        for_equal_tmp_5 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0000101"));
        for_equal_tmp_6 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0000110"));
        for_equal_tmp_7 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0000111"));
        for_equal_tmp_9 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0001001"));
        for_equal_tmp_10 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0001010"));
        for_equal_tmp_11 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0001011"));
        for_equal_tmp_12 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0001100"));
        for_equal_tmp_13 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0001101"));
        for_equal_tmp_14 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0001110"));
        for_equal_tmp_15 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0001111"));
        for_equal_tmp_17 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0010001"));
        for_equal_tmp_18 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0010010"));
        for_equal_tmp_19 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0010011"));
        for_equal_tmp_20 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0010100"));
        for_equal_tmp_21 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0010101"));
        for_equal_tmp_22 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0010110"));
        for_equal_tmp_23 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0010111"));
        for_equal_tmp_24 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0011000"));
        for_equal_tmp_25 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0011001"));
        for_equal_tmp_26 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0011010"));
        for_equal_tmp_27 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0011011"));
        for_equal_tmp_28 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0011100"));
        for_equal_tmp_29 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0011101"));
        for_equal_tmp_30 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0011110"));
        for_equal_tmp_31 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0011111"));
        for_equal_tmp_33 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0100001"));
        for_equal_tmp_34 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0100010"));
        for_equal_tmp_35 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0100011"));
        for_equal_tmp_36 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0100100"));
        for_equal_tmp_37 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0100101"));
        for_equal_tmp_38 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0100110"));
        for_equal_tmp_39 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0100111"));
        for_equal_tmp_40 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0101000"));
        for_equal_tmp_41 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0101001"));
        for_equal_tmp_42 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0101010"));
        for_equal_tmp_43 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0101011"));
        for_equal_tmp_44 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0101100"));
        for_equal_tmp_45 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0101101"));
        for_equal_tmp_46 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0101110"));
        for_equal_tmp_47 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0101111"));
        for_equal_tmp_48 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0110000"));
        for_equal_tmp_49 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0110001"));
        for_equal_tmp_50 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0110010"));
        for_equal_tmp_51 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0110011"));
        for_equal_tmp_52 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0110100"));
        for_equal_tmp_53 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0110101"));
        for_equal_tmp_54 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0110110"));
        for_equal_tmp_55 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0110111"));
        for_equal_tmp_56 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0111000"));
        for_equal_tmp_57 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0111001"));
        for_equal_tmp_58 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0111010"));
        for_equal_tmp_59 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0111011"));
        for_equal_tmp_60 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0111100"));
        for_equal_tmp_61 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0111101"));
        for_equal_tmp_62 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0111110"));
        for_equal_tmp_63 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("0111111"));
        for_equal_tmp_65 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1000001"));
        for_equal_tmp_66 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1000010"));
        for_equal_tmp_67 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1000011"));
        for_equal_tmp_68 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1000100"));
        for_equal_tmp_69 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1000101"));
        for_equal_tmp_70 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1000110"));
        for_equal_tmp_71 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1000111"));
        for_equal_tmp_72 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1001000"));
        for_equal_tmp_73 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1001001"));
        for_equal_tmp_74 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1001010"));
        for_equal_tmp_75 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1001011"));
        for_equal_tmp_76 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1001100"));
        for_equal_tmp_77 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1001101"));
        for_equal_tmp_78 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1001110"));
        for_equal_tmp_79 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1001111"));
        for_equal_tmp_80 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1010000"));
        for_equal_tmp_81 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1010001"));
        for_equal_tmp_82 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1010010"));
        for_equal_tmp_83 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1010011"));
        for_equal_tmp_84 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1010100"));
        for_equal_tmp_85 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1010101"));
        for_equal_tmp_86 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1010110"));
        for_equal_tmp_87 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1010111"));
        for_equal_tmp_88 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1011000"));
        for_equal_tmp_89 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1011001"));
        for_equal_tmp_90 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1011010"));
        for_equal_tmp_91 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1011011"));
        for_equal_tmp_92 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1011100"));
        for_equal_tmp_93 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1011101"));
        for_equal_tmp_94 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1011110"));
        for_equal_tmp_95 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1011111"));
        for_equal_tmp_96 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1100000"));
        for_equal_tmp_97 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1100001"));
        for_equal_tmp_98 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1100010"));
        for_equal_tmp_99 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1100011"));
        for_equal_tmp_100 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1100100"));
        for_equal_tmp_101 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1100101"));
        for_equal_tmp_102 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1100110"));
        for_equal_tmp_103 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1100111"));
        for_equal_tmp_104 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1101000"));
        for_equal_tmp_105 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1101001"));
        for_equal_tmp_106 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1101010"));
        for_equal_tmp_107 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1101011"));
        for_equal_tmp_108 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1101100"));
        for_equal_tmp_109 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1101101"));
        for_equal_tmp_110 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1101110"));
        for_equal_tmp_111 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1101111"));
        for_equal_tmp_112 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1110000"));
        for_equal_tmp_113 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1110001"));
        for_equal_tmp_114 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1110010"));
        for_equal_tmp_115 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1110011"));
        for_equal_tmp_116 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1110100"));
        for_equal_tmp_117 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1110101"));
        for_equal_tmp_118 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1110110"));
        for_equal_tmp_119 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1110111"));
        for_equal_tmp_120 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1111000"));
        for_equal_tmp_121 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1111001"));
        for_equal_tmp_122 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1111010"));
        for_equal_tmp_123 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1111011"));
        for_equal_tmp_124 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1111100"));
        for_equal_tmp_125 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1111101"));
        for_equal_tmp_126 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1111110"));
        for_equal_tmp_127 <= CONV_SL_1_1(i_7_0_sva_6_0=STD_LOGIC_VECTOR'("1111111"));
        for_nor_62_itm <= NOT(CONV_SL_1_1(i_7_0_sva_6_0(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000000")));
        for_nor_31_itm <= NOT((i_7_0_sva_6_0(6)) OR (i_7_0_sva_6_0(4)) OR (i_7_0_sva_6_0(3))
            OR (i_7_0_sva_6_0(2)) OR (i_7_0_sva_6_0(1)) OR (i_7_0_sva_6_0(0)));
        for_nor_15_itm <= NOT((i_7_0_sva_6_0(6)) OR (i_7_0_sva_6_0(5)) OR (i_7_0_sva_6_0(3))
            OR (i_7_0_sva_6_0(2)) OR (i_7_0_sva_6_0(1)) OR (i_7_0_sva_6_0(0)));
        for_nor_7_itm <= NOT((i_7_0_sva_6_0(6)) OR (i_7_0_sva_6_0(5)) OR (i_7_0_sva_6_0(4))
            OR (i_7_0_sva_6_0(2)) OR (i_7_0_sva_6_0(1)) OR (i_7_0_sva_6_0(0)));
        for_nor_3_itm <= NOT((i_7_0_sva_6_0(6)) OR (i_7_0_sva_6_0(5)) OR (i_7_0_sva_6_0(4))
            OR (i_7_0_sva_6_0(3)) OR (i_7_0_sva_6_0(1)) OR (i_7_0_sva_6_0(0)));
        for_nor_1_itm <= NOT((i_7_0_sva_6_0(6)) OR (i_7_0_sva_6_0(5)) OR (i_7_0_sva_6_0(4))
            OR (i_7_0_sva_6_0(3)) OR (i_7_0_sva_6_0(2)) OR (i_7_0_sva_6_0(0)));
        for_nor_itm <= NOT(CONV_SL_1_1(i_7_0_sva_6_0(6 DOWNTO 1)/=STD_LOGIC_VECTOR'("000000")));
        for_mux_itm <= MUX_v_32_128_2((input_rsci_idat(31 DOWNTO 0)), (input_rsci_idat(63
            DOWNTO 32)), (input_rsci_idat(95 DOWNTO 64)), (input_rsci_idat(127 DOWNTO
            96)), (input_rsci_idat(159 DOWNTO 128)), (input_rsci_idat(191 DOWNTO
            160)), (input_rsci_idat(223 DOWNTO 192)), (input_rsci_idat(255 DOWNTO
            224)), (input_rsci_idat(287 DOWNTO 256)), (input_rsci_idat(319 DOWNTO
            288)), (input_rsci_idat(351 DOWNTO 320)), (input_rsci_idat(383 DOWNTO
            352)), (input_rsci_idat(415 DOWNTO 384)), (input_rsci_idat(447 DOWNTO
            416)), (input_rsci_idat(479 DOWNTO 448)), (input_rsci_idat(511 DOWNTO
            480)), (input_rsci_idat(543 DOWNTO 512)), (input_rsci_idat(575 DOWNTO
            544)), (input_rsci_idat(607 DOWNTO 576)), (input_rsci_idat(639 DOWNTO
            608)), (input_rsci_idat(671 DOWNTO 640)), (input_rsci_idat(703 DOWNTO
            672)), (input_rsci_idat(735 DOWNTO 704)), (input_rsci_idat(767 DOWNTO
            736)), (input_rsci_idat(799 DOWNTO 768)), (input_rsci_idat(831 DOWNTO
            800)), (input_rsci_idat(863 DOWNTO 832)), (input_rsci_idat(895 DOWNTO
            864)), (input_rsci_idat(927 DOWNTO 896)), (input_rsci_idat(959 DOWNTO
            928)), (input_rsci_idat(991 DOWNTO 960)), (input_rsci_idat(1023 DOWNTO
            992)), (input_rsci_idat(1055 DOWNTO 1024)), (input_rsci_idat(1087 DOWNTO
            1056)), (input_rsci_idat(1119 DOWNTO 1088)), (input_rsci_idat(1151 DOWNTO
            1120)), (input_rsci_idat(1183 DOWNTO 1152)), (input_rsci_idat(1215 DOWNTO
            1184)), (input_rsci_idat(1247 DOWNTO 1216)), (input_rsci_idat(1279 DOWNTO
            1248)), (input_rsci_idat(1311 DOWNTO 1280)), (input_rsci_idat(1343 DOWNTO
            1312)), (input_rsci_idat(1375 DOWNTO 1344)), (input_rsci_idat(1407 DOWNTO
            1376)), (input_rsci_idat(1439 DOWNTO 1408)), (input_rsci_idat(1471 DOWNTO
            1440)), (input_rsci_idat(1503 DOWNTO 1472)), (input_rsci_idat(1535 DOWNTO
            1504)), (input_rsci_idat(1567 DOWNTO 1536)), (input_rsci_idat(1599 DOWNTO
            1568)), (input_rsci_idat(1631 DOWNTO 1600)), (input_rsci_idat(1663 DOWNTO
            1632)), (input_rsci_idat(1695 DOWNTO 1664)), (input_rsci_idat(1727 DOWNTO
            1696)), (input_rsci_idat(1759 DOWNTO 1728)), (input_rsci_idat(1791 DOWNTO
            1760)), (input_rsci_idat(1823 DOWNTO 1792)), (input_rsci_idat(1855 DOWNTO
            1824)), (input_rsci_idat(1887 DOWNTO 1856)), (input_rsci_idat(1919 DOWNTO
            1888)), (input_rsci_idat(1951 DOWNTO 1920)), (input_rsci_idat(1983 DOWNTO
            1952)), (input_rsci_idat(2015 DOWNTO 1984)), (input_rsci_idat(2047 DOWNTO
            2016)), (input_rsci_idat(2079 DOWNTO 2048)), (input_rsci_idat(2111 DOWNTO
            2080)), (input_rsci_idat(2143 DOWNTO 2112)), (input_rsci_idat(2175 DOWNTO
            2144)), (input_rsci_idat(2207 DOWNTO 2176)), (input_rsci_idat(2239 DOWNTO
            2208)), (input_rsci_idat(2271 DOWNTO 2240)), (input_rsci_idat(2303 DOWNTO
            2272)), (input_rsci_idat(2335 DOWNTO 2304)), (input_rsci_idat(2367 DOWNTO
            2336)), (input_rsci_idat(2399 DOWNTO 2368)), (input_rsci_idat(2431 DOWNTO
            2400)), (input_rsci_idat(2463 DOWNTO 2432)), (input_rsci_idat(2495 DOWNTO
            2464)), (input_rsci_idat(2527 DOWNTO 2496)), (input_rsci_idat(2559 DOWNTO
            2528)), (input_rsci_idat(2591 DOWNTO 2560)), (input_rsci_idat(2623 DOWNTO
            2592)), (input_rsci_idat(2655 DOWNTO 2624)), (input_rsci_idat(2687 DOWNTO
            2656)), (input_rsci_idat(2719 DOWNTO 2688)), (input_rsci_idat(2751 DOWNTO
            2720)), (input_rsci_idat(2783 DOWNTO 2752)), (input_rsci_idat(2815 DOWNTO
            2784)), (input_rsci_idat(2847 DOWNTO 2816)), (input_rsci_idat(2879 DOWNTO
            2848)), (input_rsci_idat(2911 DOWNTO 2880)), (input_rsci_idat(2943 DOWNTO
            2912)), (input_rsci_idat(2975 DOWNTO 2944)), (input_rsci_idat(3007 DOWNTO
            2976)), (input_rsci_idat(3039 DOWNTO 3008)), (input_rsci_idat(3071 DOWNTO
            3040)), (input_rsci_idat(3103 DOWNTO 3072)), (input_rsci_idat(3135 DOWNTO
            3104)), (input_rsci_idat(3167 DOWNTO 3136)), (input_rsci_idat(3199 DOWNTO
            3168)), (input_rsci_idat(3231 DOWNTO 3200)), (input_rsci_idat(3263 DOWNTO
            3232)), (input_rsci_idat(3295 DOWNTO 3264)), (input_rsci_idat(3327 DOWNTO
            3296)), (input_rsci_idat(3359 DOWNTO 3328)), (input_rsci_idat(3391 DOWNTO
            3360)), (input_rsci_idat(3423 DOWNTO 3392)), (input_rsci_idat(3455 DOWNTO
            3424)), (input_rsci_idat(3487 DOWNTO 3456)), (input_rsci_idat(3519 DOWNTO
            3488)), (input_rsci_idat(3551 DOWNTO 3520)), (input_rsci_idat(3583 DOWNTO
            3552)), (input_rsci_idat(3615 DOWNTO 3584)), (input_rsci_idat(3647 DOWNTO
            3616)), (input_rsci_idat(3679 DOWNTO 3648)), (input_rsci_idat(3711 DOWNTO
            3680)), (input_rsci_idat(3743 DOWNTO 3712)), (input_rsci_idat(3775 DOWNTO
            3744)), (input_rsci_idat(3807 DOWNTO 3776)), (input_rsci_idat(3839 DOWNTO
            3808)), (input_rsci_idat(3871 DOWNTO 3840)), (input_rsci_idat(3903 DOWNTO
            3872)), (input_rsci_idat(3935 DOWNTO 3904)), (input_rsci_idat(3967 DOWNTO
            3936)), (input_rsci_idat(3999 DOWNTO 3968)), (input_rsci_idat(4031 DOWNTO
            4000)), (input_rsci_idat(4063 DOWNTO 4032)), (input_rsci_idat(4095 DOWNTO
            4064)), i_7_0_sva_6_0);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_2047_2016_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_2047_2016_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2047_2016_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_253_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_2079_2048_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_2079_2048_lpi_2_dfm <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1,
            output_rsc_1_2079_2048_lpi_2, for_and_251_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_2015_1984_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_2015_1984_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2015_1984_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_249_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_2111_2080_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_2111_2080_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2111_2080_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_247_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_1983_1952_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_1983_1952_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1983_1952_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_245_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_2143_2112_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_2143_2112_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2143_2112_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_243_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_1951_1920_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_1951_1920_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1951_1920_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_241_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_2175_2144_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_2175_2144_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2175_2144_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_239_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_1919_1888_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_1919_1888_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1919_1888_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_237_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_2207_2176_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_2207_2176_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2207_2176_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_235_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_1887_1856_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_1887_1856_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1887_1856_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_233_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_2239_2208_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_2239_2208_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2239_2208_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_231_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_1855_1824_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_1855_1824_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1855_1824_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_229_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_2271_2240_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_2271_2240_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2271_2240_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_227_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_1823_1792_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_1823_1792_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1823_1792_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_225_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_2303_2272_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_2303_2272_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2303_2272_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_223_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_1791_1760_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_1791_1760_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1791_1760_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_221_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_2335_2304_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_2335_2304_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2335_2304_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_219_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_1759_1728_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_1759_1728_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1759_1728_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_217_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_2367_2336_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_2367_2336_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2367_2336_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_215_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_1727_1696_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_1727_1696_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1727_1696_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_213_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_2399_2368_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_2399_2368_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2399_2368_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_211_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_1695_1664_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_1695_1664_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1695_1664_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_209_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_2431_2400_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_2431_2400_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2431_2400_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_207_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_1663_1632_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_1663_1632_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1663_1632_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_205_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_2463_2432_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_2463_2432_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2463_2432_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_203_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_1631_1600_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_1631_1600_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1631_1600_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_201_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_2495_2464_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_2495_2464_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2495_2464_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_199_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_1599_1568_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_1599_1568_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1599_1568_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_197_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_2527_2496_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_2527_2496_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2527_2496_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_195_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_1567_1536_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_1567_1536_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1567_1536_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_193_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_2559_2528_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_2559_2528_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2559_2528_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_191_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_1535_1504_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_1535_1504_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1535_1504_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_189_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_2591_2560_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_2591_2560_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2591_2560_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_187_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_1503_1472_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_1503_1472_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1503_1472_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_185_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_2623_2592_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_2623_2592_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2623_2592_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_183_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_1471_1440_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_1471_1440_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1471_1440_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_181_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_2655_2624_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_2655_2624_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2655_2624_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_179_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_1439_1408_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_1439_1408_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1439_1408_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_177_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_2687_2656_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_2687_2656_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2687_2656_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_175_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_1407_1376_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_1407_1376_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1407_1376_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_173_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_2719_2688_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_2719_2688_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2719_2688_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_171_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_1375_1344_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_1375_1344_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1375_1344_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_169_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_2751_2720_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_2751_2720_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2751_2720_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_167_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_1343_1312_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_1343_1312_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1343_1312_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_165_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_2783_2752_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_2783_2752_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2783_2752_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_163_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_1311_1280_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_1311_1280_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1311_1280_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_161_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_2815_2784_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_2815_2784_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2815_2784_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_159_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_1279_1248_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_1279_1248_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1279_1248_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_157_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_2847_2816_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_2847_2816_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2847_2816_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_155_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_1247_1216_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_1247_1216_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1247_1216_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_153_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_2879_2848_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_2879_2848_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2879_2848_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_151_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_1215_1184_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_1215_1184_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1215_1184_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_149_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_2911_2880_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_2911_2880_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2911_2880_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_147_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_1183_1152_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_1183_1152_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1183_1152_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_145_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_2943_2912_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_2943_2912_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2943_2912_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_143_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_1151_1120_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_1151_1120_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1151_1120_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_141_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_2975_2944_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_2975_2944_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2975_2944_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_139_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_1119_1088_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_1119_1088_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1119_1088_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_137_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_3007_2976_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_3007_2976_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3007_2976_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_135_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_1087_1056_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_1087_1056_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1087_1056_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_133_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_3039_3008_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_3039_3008_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3039_3008_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_131_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_1055_1024_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_1055_1024_lpi_2_dfm <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1,
            output_rsc_1_1055_1024_lpi_2, for_and_129_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_3071_3040_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_3071_3040_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3071_3040_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_127_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_1023_992_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_1023_992_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1023_992_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_125_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_3103_3072_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_3103_3072_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3103_3072_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_123_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_991_960_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_991_960_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_991_960_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_121_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_3135_3104_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_3135_3104_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3135_3104_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_119_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_959_928_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_959_928_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_959_928_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_117_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_3167_3136_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_3167_3136_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3167_3136_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_115_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_927_896_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_927_896_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_927_896_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_113_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_3199_3168_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_3199_3168_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3199_3168_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_111_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_895_864_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_895_864_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_895_864_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_109_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_3231_3200_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_3231_3200_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3231_3200_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_107_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_863_832_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_863_832_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_863_832_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_105_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_3263_3232_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_3263_3232_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3263_3232_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_103_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_831_800_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_831_800_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_831_800_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_101_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_3295_3264_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_3295_3264_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3295_3264_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_99_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_799_768_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_799_768_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_799_768_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_97_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_3327_3296_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_3327_3296_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3327_3296_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_95_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_767_736_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_767_736_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_767_736_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_93_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_3359_3328_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_3359_3328_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3359_3328_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_91_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_735_704_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_735_704_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_735_704_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_89_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_3391_3360_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_3391_3360_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3391_3360_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_87_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_703_672_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_703_672_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_703_672_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_85_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_3423_3392_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_3423_3392_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3423_3392_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_83_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_671_640_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_671_640_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_671_640_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_81_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_3455_3424_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_3455_3424_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3455_3424_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_79_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_639_608_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_639_608_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_639_608_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_77_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_3487_3456_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_3487_3456_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3487_3456_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_75_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_607_576_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_607_576_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_607_576_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_73_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_3519_3488_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_3519_3488_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3519_3488_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_71_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_575_544_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_575_544_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_575_544_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_69_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_3551_3520_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_3551_3520_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3551_3520_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_67_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_543_512_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_543_512_lpi_2_dfm <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1,
            output_rsc_1_543_512_lpi_2, for_and_65_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_3583_3552_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_3583_3552_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3583_3552_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_63_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_511_480_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_511_480_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_511_480_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_61_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_3615_3584_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_3615_3584_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3615_3584_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_59_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_479_448_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_479_448_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_479_448_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_57_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_3647_3616_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_3647_3616_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3647_3616_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_55_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_447_416_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_447_416_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_447_416_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_53_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_3679_3648_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_3679_3648_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3679_3648_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_51_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_415_384_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_415_384_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_415_384_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_49_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_3711_3680_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_3711_3680_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3711_3680_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_47_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_383_352_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_383_352_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_383_352_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_45_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_3743_3712_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_3743_3712_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3743_3712_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_43_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_351_320_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_351_320_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_351_320_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_41_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_3775_3744_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_3775_3744_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3775_3744_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_39_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_319_288_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_319_288_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_319_288_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_37_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_3807_3776_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_3807_3776_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3807_3776_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_35_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_287_256_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_287_256_lpi_2_dfm <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1,
            output_rsc_1_287_256_lpi_2, for_and_33_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_3839_3808_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_3839_3808_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3839_3808_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_31_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_255_224_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_255_224_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_255_224_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_29_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_3871_3840_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_3871_3840_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3871_3840_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_27_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_223_192_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_223_192_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_223_192_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_25_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_3903_3872_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_3903_3872_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3903_3872_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_23_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_191_160_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_191_160_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_191_160_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_21_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_3935_3904_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_3935_3904_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3935_3904_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_19_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_159_128_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_159_128_lpi_2_dfm <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1,
            output_rsc_1_159_128_lpi_2, for_and_17_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_3967_3936_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_3967_3936_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3967_3936_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_15_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_127_96_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_127_96_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_127_96_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_13_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_3999_3968_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_3999_3968_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3999_3968_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_11_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_95_64_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_95_64_lpi_2_dfm <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1,
            output_rsc_1_95_64_lpi_2, for_and_9_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_4031_4000_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_4031_4000_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_4031_4000_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_7_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_63_32_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_63_32_lpi_2_dfm <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1,
            output_rsc_1_63_32_lpi_2, for_and_5_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_4063_4032_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_4063_4032_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_4063_4032_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_3_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_31_0_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_31_0_lpi_2_dfm <= output_output_mux_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_io_read_output_rsc_sdt_4095_4064_lpi_2_dfm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
      ELSIF ( or_tmp_643 = '0' ) THEN
        for_io_read_output_rsc_sdt_4095_4064_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_4095_4064_lpi_2,
            for_for_mul_1_cmx_sva_1, for_and_1_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        i_7_0_sva_1 <= STD_LOGIC_VECTOR'( "00000000");
      ELSIF ( (fsm_output(1)) = '1' ) THEN
        i_7_0_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(CONV_SIGNED(CONV_UNSIGNED(UNSIGNED(i_7_0_sva_6_0),
            7), 8) + SIGNED'( "00000001"), 8));
      END IF;
    END IF;
  END PROCESS;
  and_660_nl <= or_dcpl_330 AND (fsm_output(2));
  and_666_nl <= or_dcpl_331 AND (fsm_output(2));
  and_672_nl <= (NOT for_equal_tmp_3) AND (fsm_output(2));
  and_678_nl <= or_dcpl_332 AND (fsm_output(2));
  and_684_nl <= (NOT for_equal_tmp_5) AND (fsm_output(2));
  and_690_nl <= (NOT for_equal_tmp_6) AND (fsm_output(2));
  and_696_nl <= (NOT for_equal_tmp_7) AND (fsm_output(2));
  and_702_nl <= or_dcpl_333 AND (fsm_output(2));
  and_708_nl <= (NOT for_equal_tmp_9) AND (fsm_output(2));
  and_714_nl <= (NOT for_equal_tmp_10) AND (fsm_output(2));
  and_720_nl <= (NOT for_equal_tmp_11) AND (fsm_output(2));
  and_726_nl <= (NOT for_equal_tmp_12) AND (fsm_output(2));
  and_732_nl <= (NOT for_equal_tmp_13) AND (fsm_output(2));
  and_738_nl <= (NOT for_equal_tmp_14) AND (fsm_output(2));
  and_744_nl <= (NOT for_equal_tmp_15) AND (fsm_output(2));
  and_750_nl <= or_dcpl_334 AND (fsm_output(2));
  and_756_nl <= (NOT for_equal_tmp_17) AND (fsm_output(2));
  and_762_nl <= (NOT for_equal_tmp_18) AND (fsm_output(2));
  and_768_nl <= (NOT for_equal_tmp_19) AND (fsm_output(2));
  and_774_nl <= (NOT for_equal_tmp_20) AND (fsm_output(2));
  and_780_nl <= (NOT for_equal_tmp_21) AND (fsm_output(2));
  and_786_nl <= (NOT for_equal_tmp_22) AND (fsm_output(2));
  and_792_nl <= (NOT for_equal_tmp_23) AND (fsm_output(2));
  and_798_nl <= (NOT for_equal_tmp_24) AND (fsm_output(2));
  and_804_nl <= (NOT for_equal_tmp_25) AND (fsm_output(2));
  and_810_nl <= (NOT for_equal_tmp_26) AND (fsm_output(2));
  and_816_nl <= (NOT for_equal_tmp_27) AND (fsm_output(2));
  and_822_nl <= (NOT for_equal_tmp_28) AND (fsm_output(2));
  and_828_nl <= (NOT for_equal_tmp_29) AND (fsm_output(2));
  and_834_nl <= (NOT for_equal_tmp_30) AND (fsm_output(2));
  and_840_nl <= (NOT for_equal_tmp_31) AND (fsm_output(2));
  and_846_nl <= or_dcpl_335 AND (fsm_output(2));
  and_852_nl <= (NOT for_equal_tmp_33) AND (fsm_output(2));
  and_858_nl <= (NOT for_equal_tmp_34) AND (fsm_output(2));
  and_864_nl <= (NOT for_equal_tmp_35) AND (fsm_output(2));
  and_870_nl <= (NOT for_equal_tmp_36) AND (fsm_output(2));
  and_876_nl <= (NOT for_equal_tmp_37) AND (fsm_output(2));
  and_882_nl <= (NOT for_equal_tmp_38) AND (fsm_output(2));
  and_888_nl <= (NOT for_equal_tmp_39) AND (fsm_output(2));
  and_894_nl <= (NOT for_equal_tmp_40) AND (fsm_output(2));
  and_900_nl <= (NOT for_equal_tmp_41) AND (fsm_output(2));
  and_906_nl <= (NOT for_equal_tmp_42) AND (fsm_output(2));
  and_912_nl <= (NOT for_equal_tmp_43) AND (fsm_output(2));
  and_918_nl <= (NOT for_equal_tmp_44) AND (fsm_output(2));
  and_924_nl <= (NOT for_equal_tmp_45) AND (fsm_output(2));
  and_930_nl <= (NOT for_equal_tmp_46) AND (fsm_output(2));
  and_936_nl <= (NOT for_equal_tmp_47) AND (fsm_output(2));
  and_942_nl <= (NOT for_equal_tmp_48) AND (fsm_output(2));
  and_948_nl <= (NOT for_equal_tmp_49) AND (fsm_output(2));
  and_954_nl <= (NOT for_equal_tmp_50) AND (fsm_output(2));
  and_960_nl <= (NOT for_equal_tmp_51) AND (fsm_output(2));
  and_966_nl <= (NOT for_equal_tmp_52) AND (fsm_output(2));
  and_972_nl <= (NOT for_equal_tmp_53) AND (fsm_output(2));
  and_978_nl <= (NOT for_equal_tmp_54) AND (fsm_output(2));
  and_984_nl <= (NOT for_equal_tmp_55) AND (fsm_output(2));
  and_990_nl <= (NOT for_equal_tmp_56) AND (fsm_output(2));
  and_996_nl <= (NOT for_equal_tmp_57) AND (fsm_output(2));
  and_1002_nl <= (NOT for_equal_tmp_58) AND (fsm_output(2));
  and_1008_nl <= (NOT for_equal_tmp_59) AND (fsm_output(2));
  and_1014_nl <= (NOT for_equal_tmp_60) AND (fsm_output(2));
  and_1020_nl <= (NOT for_equal_tmp_61) AND (fsm_output(2));
  and_1026_nl <= (NOT for_equal_tmp_62) AND (fsm_output(2));
  and_1032_nl <= (NOT for_equal_tmp_63) AND (fsm_output(2));
  and_1038_nl <= or_dcpl_336 AND (fsm_output(2));
  and_1044_nl <= (NOT for_equal_tmp_65) AND (fsm_output(2));
  and_1050_nl <= (NOT for_equal_tmp_66) AND (fsm_output(2));
  and_1056_nl <= (NOT for_equal_tmp_67) AND (fsm_output(2));
  and_1062_nl <= (NOT for_equal_tmp_68) AND (fsm_output(2));
  and_1068_nl <= (NOT for_equal_tmp_69) AND (fsm_output(2));
  and_1074_nl <= (NOT for_equal_tmp_70) AND (fsm_output(2));
  and_1080_nl <= (NOT for_equal_tmp_71) AND (fsm_output(2));
  and_1086_nl <= (NOT for_equal_tmp_72) AND (fsm_output(2));
  and_1092_nl <= (NOT for_equal_tmp_73) AND (fsm_output(2));
  and_1098_nl <= (NOT for_equal_tmp_74) AND (fsm_output(2));
  and_1104_nl <= (NOT for_equal_tmp_75) AND (fsm_output(2));
  and_1110_nl <= (NOT for_equal_tmp_76) AND (fsm_output(2));
  and_1116_nl <= (NOT for_equal_tmp_77) AND (fsm_output(2));
  and_1122_nl <= (NOT for_equal_tmp_78) AND (fsm_output(2));
  and_1128_nl <= (NOT for_equal_tmp_79) AND (fsm_output(2));
  and_1134_nl <= (NOT for_equal_tmp_80) AND (fsm_output(2));
  and_1140_nl <= (NOT for_equal_tmp_81) AND (fsm_output(2));
  and_1146_nl <= (NOT for_equal_tmp_82) AND (fsm_output(2));
  and_1152_nl <= (NOT for_equal_tmp_83) AND (fsm_output(2));
  and_1158_nl <= (NOT for_equal_tmp_84) AND (fsm_output(2));
  and_1164_nl <= (NOT for_equal_tmp_85) AND (fsm_output(2));
  and_1170_nl <= (NOT for_equal_tmp_86) AND (fsm_output(2));
  and_1176_nl <= (NOT for_equal_tmp_87) AND (fsm_output(2));
  and_1182_nl <= (NOT for_equal_tmp_88) AND (fsm_output(2));
  and_1188_nl <= (NOT for_equal_tmp_89) AND (fsm_output(2));
  and_1194_nl <= (NOT for_equal_tmp_90) AND (fsm_output(2));
  and_1200_nl <= (NOT for_equal_tmp_91) AND (fsm_output(2));
  and_1206_nl <= (NOT for_equal_tmp_92) AND (fsm_output(2));
  and_1212_nl <= (NOT for_equal_tmp_93) AND (fsm_output(2));
  and_1218_nl <= (NOT for_equal_tmp_94) AND (fsm_output(2));
  and_1224_nl <= (NOT for_equal_tmp_95) AND (fsm_output(2));
  and_1230_nl <= (NOT for_equal_tmp_96) AND (fsm_output(2));
  and_1236_nl <= (NOT for_equal_tmp_97) AND (fsm_output(2));
  and_1242_nl <= (NOT for_equal_tmp_98) AND (fsm_output(2));
  and_1248_nl <= (NOT for_equal_tmp_99) AND (fsm_output(2));
  and_1254_nl <= (NOT for_equal_tmp_100) AND (fsm_output(2));
  and_1260_nl <= (NOT for_equal_tmp_101) AND (fsm_output(2));
  and_1266_nl <= (NOT for_equal_tmp_102) AND (fsm_output(2));
  and_1272_nl <= (NOT for_equal_tmp_103) AND (fsm_output(2));
  and_1278_nl <= (NOT for_equal_tmp_104) AND (fsm_output(2));
  and_1284_nl <= (NOT for_equal_tmp_105) AND (fsm_output(2));
  and_1290_nl <= (NOT for_equal_tmp_106) AND (fsm_output(2));
  and_1296_nl <= (NOT for_equal_tmp_107) AND (fsm_output(2));
  and_1302_nl <= (NOT for_equal_tmp_108) AND (fsm_output(2));
  and_1308_nl <= (NOT for_equal_tmp_109) AND (fsm_output(2));
  and_1314_nl <= (NOT for_equal_tmp_110) AND (fsm_output(2));
  and_1320_nl <= (NOT for_equal_tmp_111) AND (fsm_output(2));
  and_1326_nl <= (NOT for_equal_tmp_112) AND (fsm_output(2));
  and_1332_nl <= (NOT for_equal_tmp_113) AND (fsm_output(2));
  and_1338_nl <= (NOT for_equal_tmp_114) AND (fsm_output(2));
  and_1344_nl <= (NOT for_equal_tmp_115) AND (fsm_output(2));
  and_1350_nl <= (NOT for_equal_tmp_116) AND (fsm_output(2));
  and_1356_nl <= (NOT for_equal_tmp_117) AND (fsm_output(2));
  and_1362_nl <= (NOT for_equal_tmp_118) AND (fsm_output(2));
  and_1368_nl <= (NOT for_equal_tmp_119) AND (fsm_output(2));
  and_1374_nl <= (NOT for_equal_tmp_120) AND (fsm_output(2));
  and_1380_nl <= (NOT for_equal_tmp_121) AND (fsm_output(2));
  and_1386_nl <= (NOT for_equal_tmp_122) AND (fsm_output(2));
  and_1392_nl <= (NOT for_equal_tmp_123) AND (fsm_output(2));
  and_1398_nl <= (NOT for_equal_tmp_124) AND (fsm_output(2));
  and_1404_nl <= (NOT for_equal_tmp_125) AND (fsm_output(2));
  and_1410_nl <= (NOT for_equal_tmp_126) AND (fsm_output(2));
  and_1416_nl <= (NOT for_equal_tmp_127) AND (fsm_output(2));
  for_and_253_nl <= for_equal_tmp_63 AND (NOT or_tmp_643);
  for_and_251_nl <= or_dcpl_336 AND (NOT or_tmp_643);
  for_and_249_nl <= for_equal_tmp_62 AND (NOT or_tmp_643);
  for_and_247_nl <= for_equal_tmp_65 AND (NOT or_tmp_643);
  for_and_245_nl <= for_equal_tmp_61 AND (NOT or_tmp_643);
  for_and_243_nl <= for_equal_tmp_66 AND (NOT or_tmp_643);
  for_and_241_nl <= for_equal_tmp_60 AND (NOT or_tmp_643);
  for_and_239_nl <= for_equal_tmp_67 AND (NOT or_tmp_643);
  for_and_237_nl <= for_equal_tmp_59 AND (NOT or_tmp_643);
  for_and_235_nl <= for_equal_tmp_68 AND (NOT or_tmp_643);
  for_and_233_nl <= for_equal_tmp_58 AND (NOT or_tmp_643);
  for_and_231_nl <= for_equal_tmp_69 AND (NOT or_tmp_643);
  for_and_229_nl <= for_equal_tmp_57 AND (NOT or_tmp_643);
  for_and_227_nl <= for_equal_tmp_70 AND (NOT or_tmp_643);
  for_and_225_nl <= for_equal_tmp_56 AND (NOT or_tmp_643);
  for_and_223_nl <= for_equal_tmp_71 AND (NOT or_tmp_643);
  for_and_221_nl <= for_equal_tmp_55 AND (NOT or_tmp_643);
  for_and_219_nl <= for_equal_tmp_72 AND (NOT or_tmp_643);
  for_and_217_nl <= for_equal_tmp_54 AND (NOT or_tmp_643);
  for_and_215_nl <= for_equal_tmp_73 AND (NOT or_tmp_643);
  for_and_213_nl <= for_equal_tmp_53 AND (NOT or_tmp_643);
  for_and_211_nl <= for_equal_tmp_74 AND (NOT or_tmp_643);
  for_and_209_nl <= for_equal_tmp_52 AND (NOT or_tmp_643);
  for_and_207_nl <= for_equal_tmp_75 AND (NOT or_tmp_643);
  for_and_205_nl <= for_equal_tmp_51 AND (NOT or_tmp_643);
  for_and_203_nl <= for_equal_tmp_76 AND (NOT or_tmp_643);
  for_and_201_nl <= for_equal_tmp_50 AND (NOT or_tmp_643);
  for_and_199_nl <= for_equal_tmp_77 AND (NOT or_tmp_643);
  for_and_197_nl <= for_equal_tmp_49 AND (NOT or_tmp_643);
  for_and_195_nl <= for_equal_tmp_78 AND (NOT or_tmp_643);
  for_and_193_nl <= for_equal_tmp_48 AND (NOT or_tmp_643);
  for_and_191_nl <= for_equal_tmp_79 AND (NOT or_tmp_643);
  for_and_189_nl <= for_equal_tmp_47 AND (NOT or_tmp_643);
  for_and_187_nl <= for_equal_tmp_80 AND (NOT or_tmp_643);
  for_and_185_nl <= for_equal_tmp_46 AND (NOT or_tmp_643);
  for_and_183_nl <= for_equal_tmp_81 AND (NOT or_tmp_643);
  for_and_181_nl <= for_equal_tmp_45 AND (NOT or_tmp_643);
  for_and_179_nl <= for_equal_tmp_82 AND (NOT or_tmp_643);
  for_and_177_nl <= for_equal_tmp_44 AND (NOT or_tmp_643);
  for_and_175_nl <= for_equal_tmp_83 AND (NOT or_tmp_643);
  for_and_173_nl <= for_equal_tmp_43 AND (NOT or_tmp_643);
  for_and_171_nl <= for_equal_tmp_84 AND (NOT or_tmp_643);
  for_and_169_nl <= for_equal_tmp_42 AND (NOT or_tmp_643);
  for_and_167_nl <= for_equal_tmp_85 AND (NOT or_tmp_643);
  for_and_165_nl <= for_equal_tmp_41 AND (NOT or_tmp_643);
  for_and_163_nl <= for_equal_tmp_86 AND (NOT or_tmp_643);
  for_and_161_nl <= for_equal_tmp_40 AND (NOT or_tmp_643);
  for_and_159_nl <= for_equal_tmp_87 AND (NOT or_tmp_643);
  for_and_157_nl <= for_equal_tmp_39 AND (NOT or_tmp_643);
  for_and_155_nl <= for_equal_tmp_88 AND (NOT or_tmp_643);
  for_and_153_nl <= for_equal_tmp_38 AND (NOT or_tmp_643);
  for_and_151_nl <= for_equal_tmp_89 AND (NOT or_tmp_643);
  for_and_149_nl <= for_equal_tmp_37 AND (NOT or_tmp_643);
  for_and_147_nl <= for_equal_tmp_90 AND (NOT or_tmp_643);
  for_and_145_nl <= for_equal_tmp_36 AND (NOT or_tmp_643);
  for_and_143_nl <= for_equal_tmp_91 AND (NOT or_tmp_643);
  for_and_141_nl <= for_equal_tmp_35 AND (NOT or_tmp_643);
  for_and_139_nl <= for_equal_tmp_92 AND (NOT or_tmp_643);
  for_and_137_nl <= for_equal_tmp_34 AND (NOT or_tmp_643);
  for_and_135_nl <= for_equal_tmp_93 AND (NOT or_tmp_643);
  for_and_133_nl <= for_equal_tmp_33 AND (NOT or_tmp_643);
  for_and_131_nl <= for_equal_tmp_94 AND (NOT or_tmp_643);
  for_and_129_nl <= or_dcpl_335 AND (NOT or_tmp_643);
  for_and_127_nl <= for_equal_tmp_95 AND (NOT or_tmp_643);
  for_and_125_nl <= for_equal_tmp_31 AND (NOT or_tmp_643);
  for_and_123_nl <= for_equal_tmp_96 AND (NOT or_tmp_643);
  for_and_121_nl <= for_equal_tmp_30 AND (NOT or_tmp_643);
  for_and_119_nl <= for_equal_tmp_97 AND (NOT or_tmp_643);
  for_and_117_nl <= for_equal_tmp_29 AND (NOT or_tmp_643);
  for_and_115_nl <= for_equal_tmp_98 AND (NOT or_tmp_643);
  for_and_113_nl <= for_equal_tmp_28 AND (NOT or_tmp_643);
  for_and_111_nl <= for_equal_tmp_99 AND (NOT or_tmp_643);
  for_and_109_nl <= for_equal_tmp_27 AND (NOT or_tmp_643);
  for_and_107_nl <= for_equal_tmp_100 AND (NOT or_tmp_643);
  for_and_105_nl <= for_equal_tmp_26 AND (NOT or_tmp_643);
  for_and_103_nl <= for_equal_tmp_101 AND (NOT or_tmp_643);
  for_and_101_nl <= for_equal_tmp_25 AND (NOT or_tmp_643);
  for_and_99_nl <= for_equal_tmp_102 AND (NOT or_tmp_643);
  for_and_97_nl <= for_equal_tmp_24 AND (NOT or_tmp_643);
  for_and_95_nl <= for_equal_tmp_103 AND (NOT or_tmp_643);
  for_and_93_nl <= for_equal_tmp_23 AND (NOT or_tmp_643);
  for_and_91_nl <= for_equal_tmp_104 AND (NOT or_tmp_643);
  for_and_89_nl <= for_equal_tmp_22 AND (NOT or_tmp_643);
  for_and_87_nl <= for_equal_tmp_105 AND (NOT or_tmp_643);
  for_and_85_nl <= for_equal_tmp_21 AND (NOT or_tmp_643);
  for_and_83_nl <= for_equal_tmp_106 AND (NOT or_tmp_643);
  for_and_81_nl <= for_equal_tmp_20 AND (NOT or_tmp_643);
  for_and_79_nl <= for_equal_tmp_107 AND (NOT or_tmp_643);
  for_and_77_nl <= for_equal_tmp_19 AND (NOT or_tmp_643);
  for_and_75_nl <= for_equal_tmp_108 AND (NOT or_tmp_643);
  for_and_73_nl <= for_equal_tmp_18 AND (NOT or_tmp_643);
  for_and_71_nl <= for_equal_tmp_109 AND (NOT or_tmp_643);
  for_and_69_nl <= for_equal_tmp_17 AND (NOT or_tmp_643);
  for_and_67_nl <= for_equal_tmp_110 AND (NOT or_tmp_643);
  for_and_65_nl <= or_dcpl_334 AND (NOT or_tmp_643);
  for_and_63_nl <= for_equal_tmp_111 AND (NOT or_tmp_643);
  for_and_61_nl <= for_equal_tmp_15 AND (NOT or_tmp_643);
  for_and_59_nl <= for_equal_tmp_112 AND (NOT or_tmp_643);
  for_and_57_nl <= for_equal_tmp_14 AND (NOT or_tmp_643);
  for_and_55_nl <= for_equal_tmp_113 AND (NOT or_tmp_643);
  for_and_53_nl <= for_equal_tmp_13 AND (NOT or_tmp_643);
  for_and_51_nl <= for_equal_tmp_114 AND (NOT or_tmp_643);
  for_and_49_nl <= for_equal_tmp_12 AND (NOT or_tmp_643);
  for_and_47_nl <= for_equal_tmp_115 AND (NOT or_tmp_643);
  for_and_45_nl <= for_equal_tmp_11 AND (NOT or_tmp_643);
  for_and_43_nl <= for_equal_tmp_116 AND (NOT or_tmp_643);
  for_and_41_nl <= for_equal_tmp_10 AND (NOT or_tmp_643);
  for_and_39_nl <= for_equal_tmp_117 AND (NOT or_tmp_643);
  for_and_37_nl <= for_equal_tmp_9 AND (NOT or_tmp_643);
  for_and_35_nl <= for_equal_tmp_118 AND (NOT or_tmp_643);
  for_and_33_nl <= or_dcpl_333 AND (NOT or_tmp_643);
  for_and_31_nl <= for_equal_tmp_119 AND (NOT or_tmp_643);
  for_and_29_nl <= for_equal_tmp_7 AND (NOT or_tmp_643);
  for_and_27_nl <= for_equal_tmp_120 AND (NOT or_tmp_643);
  for_and_25_nl <= for_equal_tmp_6 AND (NOT or_tmp_643);
  for_and_23_nl <= for_equal_tmp_121 AND (NOT or_tmp_643);
  for_and_21_nl <= for_equal_tmp_5 AND (NOT or_tmp_643);
  for_and_19_nl <= for_equal_tmp_122 AND (NOT or_tmp_643);
  for_and_17_nl <= or_dcpl_332 AND (NOT or_tmp_643);
  for_and_15_nl <= for_equal_tmp_123 AND (NOT or_tmp_643);
  for_and_13_nl <= for_equal_tmp_3 AND (NOT or_tmp_643);
  for_and_11_nl <= for_equal_tmp_124 AND (NOT or_tmp_643);
  for_and_9_nl <= or_dcpl_331 AND (NOT or_tmp_643);
  for_and_7_nl <= for_equal_tmp_125 AND (NOT or_tmp_643);
  for_and_5_nl <= or_dcpl_330 AND (NOT or_tmp_643);
  for_and_3_nl <= for_equal_tmp_126 AND (NOT or_tmp_643);
  for_and_1_nl <= for_equal_tmp_127 AND (NOT or_tmp_643);
END v1;

-- ------------------------------------------------------------------
--  Design Unit:    fir
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.ccs_out_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;


ENTITY fir IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    input_rsc_dat : IN STD_LOGIC_VECTOR (4095 DOWNTO 0);
    input_rsc_triosy_lz : OUT STD_LOGIC;
    output_rsc_dat : OUT STD_LOGIC_VECTOR (4095 DOWNTO 0);
    output_rsc_triosy_lz : OUT STD_LOGIC
  );
END fir;

ARCHITECTURE v1 OF fir IS
  -- Default Constants

  COMPONENT fir_core
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      input_rsc_dat : IN STD_LOGIC_VECTOR (4095 DOWNTO 0);
      input_rsc_triosy_lz : OUT STD_LOGIC;
      output_rsc_dat : OUT STD_LOGIC_VECTOR (4095 DOWNTO 0);
      output_rsc_triosy_lz : OUT STD_LOGIC
    );
  END COMPONENT;
  SIGNAL fir_core_inst_input_rsc_dat : STD_LOGIC_VECTOR (4095 DOWNTO 0);
  SIGNAL fir_core_inst_output_rsc_dat : STD_LOGIC_VECTOR (4095 DOWNTO 0);

BEGIN
  fir_core_inst : fir_core
    PORT MAP(
      clk => clk,
      rst => rst,
      input_rsc_dat => fir_core_inst_input_rsc_dat,
      input_rsc_triosy_lz => input_rsc_triosy_lz,
      output_rsc_dat => fir_core_inst_output_rsc_dat,
      output_rsc_triosy_lz => output_rsc_triosy_lz
    );
  fir_core_inst_input_rsc_dat <= input_rsc_dat;
  output_rsc_dat <= fir_core_inst_output_rsc_dat;

END v1;



