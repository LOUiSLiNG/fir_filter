
//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/ccs_out_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module ccs_out_v1 (dat, idat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output   [width-1:0] dat;
  input    [width-1:0] idat;

  wire     [width-1:0] dat;

  assign dat = idat;

endmodule




//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   dss545@hansolo.poly.edu
//  Generated date: Wed Feb  3 19:34:32 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    fir_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module fir_core_core_fsm (
  clk, rst, fsm_output, for_C_2_tr0
);
  input clk;
  input rst;
  output [4:0] fsm_output;
  reg [4:0] fsm_output;
  input for_C_2_tr0;


  // FSM State Type Declaration for fir_core_core_fsm_1
  parameter
    main_C_0 = 3'd0,
    for_C_0 = 3'd1,
    for_C_1 = 3'd2,
    for_C_2 = 3'd3,
    main_C_1 = 3'd4;

  reg [2:0] state_var;
  reg [2:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : fir_core_core_fsm_1
    case (state_var)
      for_C_0 : begin
        fsm_output = 5'b00010;
        state_var_NS = for_C_1;
      end
      for_C_1 : begin
        fsm_output = 5'b00100;
        state_var_NS = for_C_2;
      end
      for_C_2 : begin
        fsm_output = 5'b01000;
        if ( for_C_2_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = for_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 5'b10000;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 5'b00001;
        state_var_NS = for_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= main_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    fir_core
// ------------------------------------------------------------------


module fir_core (
  clk, rst, input_rsc_dat, input_rsc_triosy_lz, output_rsc_dat, output_rsc_triosy_lz
);
  input clk;
  input rst;
  input [4095:0] input_rsc_dat;
  output input_rsc_triosy_lz;
  output [4095:0] output_rsc_dat;
  output output_rsc_triosy_lz;


  // Interconnect Declarations
  wire [4095:0] input_rsci_idat;
  reg [31:0] output_rsci_idat_4095_4064;
  reg [31:0] output_rsci_idat_4063_4032;
  reg [31:0] output_rsci_idat_4031_4000;
  reg [31:0] output_rsci_idat_3999_3968;
  reg [31:0] output_rsci_idat_3967_3936;
  reg [31:0] output_rsci_idat_3935_3904;
  reg [31:0] output_rsci_idat_3903_3872;
  reg [31:0] output_rsci_idat_3871_3840;
  reg [31:0] output_rsci_idat_3839_3808;
  reg [31:0] output_rsci_idat_3807_3776;
  reg [31:0] output_rsci_idat_3775_3744;
  reg [31:0] output_rsci_idat_3743_3712;
  reg [31:0] output_rsci_idat_3711_3680;
  reg [31:0] output_rsci_idat_3679_3648;
  reg [31:0] output_rsci_idat_3647_3616;
  reg [31:0] output_rsci_idat_3615_3584;
  reg [31:0] output_rsci_idat_3583_3552;
  reg [31:0] output_rsci_idat_3551_3520;
  reg [31:0] output_rsci_idat_3519_3488;
  reg [31:0] output_rsci_idat_3487_3456;
  reg [31:0] output_rsci_idat_3455_3424;
  reg [31:0] output_rsci_idat_3423_3392;
  reg [31:0] output_rsci_idat_3391_3360;
  reg [31:0] output_rsci_idat_3359_3328;
  reg [31:0] output_rsci_idat_3327_3296;
  reg [31:0] output_rsci_idat_3295_3264;
  reg [31:0] output_rsci_idat_3263_3232;
  reg [31:0] output_rsci_idat_3231_3200;
  reg [31:0] output_rsci_idat_3199_3168;
  reg [31:0] output_rsci_idat_3167_3136;
  reg [31:0] output_rsci_idat_3135_3104;
  reg [31:0] output_rsci_idat_3103_3072;
  reg [31:0] output_rsci_idat_3071_3040;
  reg [31:0] output_rsci_idat_3039_3008;
  reg [31:0] output_rsci_idat_3007_2976;
  reg [31:0] output_rsci_idat_2975_2944;
  reg [31:0] output_rsci_idat_2943_2912;
  reg [31:0] output_rsci_idat_2911_2880;
  reg [31:0] output_rsci_idat_2879_2848;
  reg [31:0] output_rsci_idat_2847_2816;
  reg [31:0] output_rsci_idat_2815_2784;
  reg [31:0] output_rsci_idat_2783_2752;
  reg [31:0] output_rsci_idat_2751_2720;
  reg [31:0] output_rsci_idat_2719_2688;
  reg [31:0] output_rsci_idat_2687_2656;
  reg [31:0] output_rsci_idat_2655_2624;
  reg [31:0] output_rsci_idat_2623_2592;
  reg [31:0] output_rsci_idat_2591_2560;
  reg [31:0] output_rsci_idat_2559_2528;
  reg [31:0] output_rsci_idat_2527_2496;
  reg [31:0] output_rsci_idat_2495_2464;
  reg [31:0] output_rsci_idat_2463_2432;
  reg [31:0] output_rsci_idat_2431_2400;
  reg [31:0] output_rsci_idat_2399_2368;
  reg [31:0] output_rsci_idat_2367_2336;
  reg [31:0] output_rsci_idat_2335_2304;
  reg [31:0] output_rsci_idat_2303_2272;
  reg [31:0] output_rsci_idat_2271_2240;
  reg [31:0] output_rsci_idat_2239_2208;
  reg [31:0] output_rsci_idat_2207_2176;
  reg [31:0] output_rsci_idat_2175_2144;
  reg [31:0] output_rsci_idat_2143_2112;
  reg [31:0] output_rsci_idat_2111_2080;
  reg [31:0] output_rsci_idat_2079_2048;
  reg [31:0] output_rsci_idat_2047_2016;
  reg [31:0] output_rsci_idat_2015_1984;
  reg [31:0] output_rsci_idat_1983_1952;
  reg [31:0] output_rsci_idat_1951_1920;
  reg [31:0] output_rsci_idat_1919_1888;
  reg [31:0] output_rsci_idat_1887_1856;
  reg [31:0] output_rsci_idat_1855_1824;
  reg [31:0] output_rsci_idat_1823_1792;
  reg [31:0] output_rsci_idat_1791_1760;
  reg [31:0] output_rsci_idat_1759_1728;
  reg [31:0] output_rsci_idat_1727_1696;
  reg [31:0] output_rsci_idat_1695_1664;
  reg [31:0] output_rsci_idat_1663_1632;
  reg [31:0] output_rsci_idat_1631_1600;
  reg [31:0] output_rsci_idat_1599_1568;
  reg [31:0] output_rsci_idat_1567_1536;
  reg [31:0] output_rsci_idat_1535_1504;
  reg [31:0] output_rsci_idat_1503_1472;
  reg [31:0] output_rsci_idat_1471_1440;
  reg [31:0] output_rsci_idat_1439_1408;
  reg [31:0] output_rsci_idat_1407_1376;
  reg [31:0] output_rsci_idat_1375_1344;
  reg [31:0] output_rsci_idat_1343_1312;
  reg [31:0] output_rsci_idat_1311_1280;
  reg [31:0] output_rsci_idat_1279_1248;
  reg [31:0] output_rsci_idat_1247_1216;
  reg [31:0] output_rsci_idat_1215_1184;
  reg [31:0] output_rsci_idat_1183_1152;
  reg [31:0] output_rsci_idat_1151_1120;
  reg [31:0] output_rsci_idat_1119_1088;
  reg [31:0] output_rsci_idat_1087_1056;
  reg [31:0] output_rsci_idat_1055_1024;
  reg [31:0] output_rsci_idat_1023_992;
  reg [31:0] output_rsci_idat_991_960;
  reg [31:0] output_rsci_idat_959_928;
  reg [31:0] output_rsci_idat_927_896;
  reg [31:0] output_rsci_idat_895_864;
  reg [31:0] output_rsci_idat_863_832;
  reg [31:0] output_rsci_idat_831_800;
  reg [31:0] output_rsci_idat_799_768;
  reg [31:0] output_rsci_idat_767_736;
  reg [31:0] output_rsci_idat_735_704;
  reg [31:0] output_rsci_idat_703_672;
  reg [31:0] output_rsci_idat_671_640;
  reg [31:0] output_rsci_idat_639_608;
  reg [31:0] output_rsci_idat_607_576;
  reg [31:0] output_rsci_idat_575_544;
  reg [31:0] output_rsci_idat_543_512;
  reg [31:0] output_rsci_idat_511_480;
  reg [31:0] output_rsci_idat_479_448;
  reg [31:0] output_rsci_idat_447_416;
  reg [31:0] output_rsci_idat_415_384;
  reg [31:0] output_rsci_idat_383_352;
  reg [31:0] output_rsci_idat_351_320;
  reg [31:0] output_rsci_idat_319_288;
  reg [31:0] output_rsci_idat_287_256;
  reg [31:0] output_rsci_idat_255_224;
  reg [31:0] output_rsci_idat_223_192;
  reg [31:0] output_rsci_idat_191_160;
  reg [31:0] output_rsci_idat_159_128;
  reg [31:0] output_rsci_idat_127_96;
  reg [31:0] output_rsci_idat_95_64;
  reg [31:0] output_rsci_idat_63_32;
  reg [31:0] output_rsci_idat_31_0;
  wire [4:0] fsm_output;
  wire for_or_tmp;
  wire or_dcpl_330;
  wire or_dcpl_331;
  wire or_dcpl_332;
  wire or_dcpl_333;
  wire or_dcpl_334;
  wire or_dcpl_335;
  wire or_dcpl_336;
  wire or_tmp_259;
  wire or_tmp_643;
  reg for_nor_62_itm;
  reg for_nor_31_itm;
  reg for_nor_15_itm;
  reg for_nor_7_itm;
  reg for_nor_3_itm;
  reg for_nor_1_itm;
  reg for_nor_itm;
  reg [6:0] i_7_0_sva_6_0;
  reg [7:0] i_7_0_sva_1;
  wire [8:0] nl_i_7_0_sva_1;
  reg for_equal_tmp_3;
  reg for_equal_tmp_5;
  reg for_equal_tmp_6;
  reg for_equal_tmp_7;
  reg for_equal_tmp_9;
  reg for_equal_tmp_10;
  reg for_equal_tmp_11;
  reg for_equal_tmp_12;
  reg for_equal_tmp_13;
  reg for_equal_tmp_14;
  reg for_equal_tmp_15;
  reg for_equal_tmp_17;
  reg for_equal_tmp_18;
  reg for_equal_tmp_19;
  reg for_equal_tmp_20;
  reg for_equal_tmp_21;
  reg for_equal_tmp_22;
  reg for_equal_tmp_23;
  reg for_equal_tmp_24;
  reg for_equal_tmp_25;
  reg for_equal_tmp_26;
  reg for_equal_tmp_27;
  reg for_equal_tmp_28;
  reg for_equal_tmp_29;
  reg for_equal_tmp_30;
  reg for_equal_tmp_31;
  reg for_equal_tmp_33;
  reg for_equal_tmp_34;
  reg for_equal_tmp_35;
  reg for_equal_tmp_36;
  reg for_equal_tmp_37;
  reg for_equal_tmp_38;
  reg for_equal_tmp_39;
  reg for_equal_tmp_40;
  reg for_equal_tmp_41;
  reg for_equal_tmp_42;
  reg for_equal_tmp_43;
  reg for_equal_tmp_44;
  reg for_equal_tmp_45;
  reg for_equal_tmp_46;
  reg for_equal_tmp_47;
  reg for_equal_tmp_48;
  reg for_equal_tmp_49;
  reg for_equal_tmp_50;
  reg for_equal_tmp_51;
  reg for_equal_tmp_52;
  reg for_equal_tmp_53;
  reg for_equal_tmp_54;
  reg for_equal_tmp_55;
  reg for_equal_tmp_56;
  reg for_equal_tmp_57;
  reg for_equal_tmp_58;
  reg for_equal_tmp_59;
  reg for_equal_tmp_60;
  reg for_equal_tmp_61;
  reg for_equal_tmp_62;
  reg for_equal_tmp_63;
  reg for_equal_tmp_65;
  reg for_equal_tmp_66;
  reg for_equal_tmp_67;
  reg for_equal_tmp_68;
  reg for_equal_tmp_69;
  reg for_equal_tmp_70;
  reg for_equal_tmp_71;
  reg for_equal_tmp_72;
  reg for_equal_tmp_73;
  reg for_equal_tmp_74;
  reg for_equal_tmp_75;
  reg for_equal_tmp_76;
  reg for_equal_tmp_77;
  reg for_equal_tmp_78;
  reg for_equal_tmp_79;
  reg for_equal_tmp_80;
  reg for_equal_tmp_81;
  reg for_equal_tmp_82;
  reg for_equal_tmp_83;
  reg for_equal_tmp_84;
  reg for_equal_tmp_85;
  reg for_equal_tmp_86;
  reg for_equal_tmp_87;
  reg for_equal_tmp_88;
  reg for_equal_tmp_89;
  reg for_equal_tmp_90;
  reg for_equal_tmp_91;
  reg for_equal_tmp_92;
  reg for_equal_tmp_93;
  reg for_equal_tmp_94;
  reg for_equal_tmp_95;
  reg for_equal_tmp_96;
  reg for_equal_tmp_97;
  reg for_equal_tmp_98;
  reg for_equal_tmp_99;
  reg for_equal_tmp_100;
  reg for_equal_tmp_101;
  reg for_equal_tmp_102;
  reg for_equal_tmp_103;
  reg for_equal_tmp_104;
  reg for_equal_tmp_105;
  reg for_equal_tmp_106;
  reg for_equal_tmp_107;
  reg for_equal_tmp_108;
  reg for_equal_tmp_109;
  reg for_equal_tmp_110;
  reg for_equal_tmp_111;
  reg for_equal_tmp_112;
  reg for_equal_tmp_113;
  reg for_equal_tmp_114;
  reg for_equal_tmp_115;
  reg for_equal_tmp_116;
  reg for_equal_tmp_117;
  reg for_equal_tmp_118;
  reg for_equal_tmp_119;
  reg for_equal_tmp_120;
  reg for_equal_tmp_121;
  reg for_equal_tmp_122;
  reg for_equal_tmp_123;
  reg for_equal_tmp_124;
  reg for_equal_tmp_125;
  reg for_equal_tmp_126;
  reg for_equal_tmp_127;
  reg reg_output_rsc_triosy_obj_ld_cse;
  wire [31:0] output_output_mux_cse;
  reg [31:0] output_rsc_1_2047_2016_lpi_2;
  reg [31:0] output_rsc_1_2079_2048_lpi_2;
  reg [31:0] output_rsc_1_2015_1984_lpi_2;
  reg [31:0] output_rsc_1_2111_2080_lpi_2;
  reg [31:0] output_rsc_1_1983_1952_lpi_2;
  reg [31:0] output_rsc_1_2143_2112_lpi_2;
  reg [31:0] output_rsc_1_1951_1920_lpi_2;
  reg [31:0] output_rsc_1_2175_2144_lpi_2;
  reg [31:0] output_rsc_1_1919_1888_lpi_2;
  reg [31:0] output_rsc_1_2207_2176_lpi_2;
  reg [31:0] output_rsc_1_1887_1856_lpi_2;
  reg [31:0] output_rsc_1_2239_2208_lpi_2;
  reg [31:0] output_rsc_1_1855_1824_lpi_2;
  reg [31:0] output_rsc_1_2271_2240_lpi_2;
  reg [31:0] output_rsc_1_1823_1792_lpi_2;
  reg [31:0] output_rsc_1_2303_2272_lpi_2;
  reg [31:0] output_rsc_1_1791_1760_lpi_2;
  reg [31:0] output_rsc_1_2335_2304_lpi_2;
  reg [31:0] output_rsc_1_1759_1728_lpi_2;
  reg [31:0] output_rsc_1_2367_2336_lpi_2;
  reg [31:0] output_rsc_1_1727_1696_lpi_2;
  reg [31:0] output_rsc_1_2399_2368_lpi_2;
  reg [31:0] output_rsc_1_1695_1664_lpi_2;
  reg [31:0] output_rsc_1_2431_2400_lpi_2;
  reg [31:0] output_rsc_1_1663_1632_lpi_2;
  reg [31:0] output_rsc_1_2463_2432_lpi_2;
  reg [31:0] output_rsc_1_1631_1600_lpi_2;
  reg [31:0] output_rsc_1_2495_2464_lpi_2;
  reg [31:0] output_rsc_1_1599_1568_lpi_2;
  reg [31:0] output_rsc_1_2527_2496_lpi_2;
  reg [31:0] output_rsc_1_1567_1536_lpi_2;
  reg [31:0] output_rsc_1_2559_2528_lpi_2;
  reg [31:0] output_rsc_1_1535_1504_lpi_2;
  reg [31:0] output_rsc_1_2591_2560_lpi_2;
  reg [31:0] output_rsc_1_1503_1472_lpi_2;
  reg [31:0] output_rsc_1_2623_2592_lpi_2;
  reg [31:0] output_rsc_1_1471_1440_lpi_2;
  reg [31:0] output_rsc_1_2655_2624_lpi_2;
  reg [31:0] output_rsc_1_1439_1408_lpi_2;
  reg [31:0] output_rsc_1_2687_2656_lpi_2;
  reg [31:0] output_rsc_1_1407_1376_lpi_2;
  reg [31:0] output_rsc_1_2719_2688_lpi_2;
  reg [31:0] output_rsc_1_1375_1344_lpi_2;
  reg [31:0] output_rsc_1_2751_2720_lpi_2;
  reg [31:0] output_rsc_1_1343_1312_lpi_2;
  reg [31:0] output_rsc_1_2783_2752_lpi_2;
  reg [31:0] output_rsc_1_1311_1280_lpi_2;
  reg [31:0] output_rsc_1_2815_2784_lpi_2;
  reg [31:0] output_rsc_1_1279_1248_lpi_2;
  reg [31:0] output_rsc_1_2847_2816_lpi_2;
  reg [31:0] output_rsc_1_1247_1216_lpi_2;
  reg [31:0] output_rsc_1_2879_2848_lpi_2;
  reg [31:0] output_rsc_1_1215_1184_lpi_2;
  reg [31:0] output_rsc_1_2911_2880_lpi_2;
  reg [31:0] output_rsc_1_1183_1152_lpi_2;
  reg [31:0] output_rsc_1_2943_2912_lpi_2;
  reg [31:0] output_rsc_1_1151_1120_lpi_2;
  reg [31:0] output_rsc_1_2975_2944_lpi_2;
  reg [31:0] output_rsc_1_1119_1088_lpi_2;
  reg [31:0] output_rsc_1_3007_2976_lpi_2;
  reg [31:0] output_rsc_1_1087_1056_lpi_2;
  reg [31:0] output_rsc_1_3039_3008_lpi_2;
  reg [31:0] output_rsc_1_1055_1024_lpi_2;
  reg [31:0] output_rsc_1_3071_3040_lpi_2;
  reg [31:0] output_rsc_1_1023_992_lpi_2;
  reg [31:0] output_rsc_1_3103_3072_lpi_2;
  reg [31:0] output_rsc_1_991_960_lpi_2;
  reg [31:0] output_rsc_1_3135_3104_lpi_2;
  reg [31:0] output_rsc_1_959_928_lpi_2;
  reg [31:0] output_rsc_1_3167_3136_lpi_2;
  reg [31:0] output_rsc_1_927_896_lpi_2;
  reg [31:0] output_rsc_1_3199_3168_lpi_2;
  reg [31:0] output_rsc_1_895_864_lpi_2;
  reg [31:0] output_rsc_1_3231_3200_lpi_2;
  reg [31:0] output_rsc_1_863_832_lpi_2;
  reg [31:0] output_rsc_1_3263_3232_lpi_2;
  reg [31:0] output_rsc_1_831_800_lpi_2;
  reg [31:0] output_rsc_1_3295_3264_lpi_2;
  reg [31:0] output_rsc_1_799_768_lpi_2;
  reg [31:0] output_rsc_1_3327_3296_lpi_2;
  reg [31:0] output_rsc_1_767_736_lpi_2;
  reg [31:0] output_rsc_1_3359_3328_lpi_2;
  reg [31:0] output_rsc_1_735_704_lpi_2;
  reg [31:0] output_rsc_1_3391_3360_lpi_2;
  reg [31:0] output_rsc_1_703_672_lpi_2;
  reg [31:0] output_rsc_1_3423_3392_lpi_2;
  reg [31:0] output_rsc_1_671_640_lpi_2;
  reg [31:0] output_rsc_1_3455_3424_lpi_2;
  reg [31:0] output_rsc_1_639_608_lpi_2;
  reg [31:0] output_rsc_1_3487_3456_lpi_2;
  reg [31:0] output_rsc_1_607_576_lpi_2;
  reg [31:0] output_rsc_1_3519_3488_lpi_2;
  reg [31:0] output_rsc_1_575_544_lpi_2;
  reg [31:0] output_rsc_1_3551_3520_lpi_2;
  reg [31:0] output_rsc_1_543_512_lpi_2;
  reg [31:0] output_rsc_1_3583_3552_lpi_2;
  reg [31:0] output_rsc_1_511_480_lpi_2;
  reg [31:0] output_rsc_1_3615_3584_lpi_2;
  reg [31:0] output_rsc_1_479_448_lpi_2;
  reg [31:0] output_rsc_1_3647_3616_lpi_2;
  reg [31:0] output_rsc_1_447_416_lpi_2;
  reg [31:0] output_rsc_1_3679_3648_lpi_2;
  reg [31:0] output_rsc_1_415_384_lpi_2;
  reg [31:0] output_rsc_1_3711_3680_lpi_2;
  reg [31:0] output_rsc_1_383_352_lpi_2;
  reg [31:0] output_rsc_1_3743_3712_lpi_2;
  reg [31:0] output_rsc_1_351_320_lpi_2;
  reg [31:0] output_rsc_1_3775_3744_lpi_2;
  reg [31:0] output_rsc_1_319_288_lpi_2;
  reg [31:0] output_rsc_1_3807_3776_lpi_2;
  reg [31:0] output_rsc_1_287_256_lpi_2;
  reg [31:0] output_rsc_1_3839_3808_lpi_2;
  reg [31:0] output_rsc_1_255_224_lpi_2;
  reg [31:0] output_rsc_1_3871_3840_lpi_2;
  reg [31:0] output_rsc_1_223_192_lpi_2;
  reg [31:0] output_rsc_1_3903_3872_lpi_2;
  reg [31:0] output_rsc_1_191_160_lpi_2;
  reg [31:0] output_rsc_1_3935_3904_lpi_2;
  reg [31:0] output_rsc_1_159_128_lpi_2;
  reg [31:0] output_rsc_1_3967_3936_lpi_2;
  reg [31:0] output_rsc_1_127_96_lpi_2;
  reg [31:0] output_rsc_1_3999_3968_lpi_2;
  reg [31:0] output_rsc_1_95_64_lpi_2;
  reg [31:0] output_rsc_1_4031_4000_lpi_2;
  reg [31:0] output_rsc_1_63_32_lpi_2;
  reg [31:0] output_rsc_1_4063_4032_lpi_2;
  reg [31:0] output_rsc_1_31_0_lpi_2;
  reg [31:0] output_rsc_1_4095_4064_lpi_2;
  reg [31:0] for_io_read_output_rsc_sdt_4095_4064_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_4063_4032_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_4031_4000_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_3999_3968_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_3967_3936_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_3935_3904_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_3903_3872_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_3871_3840_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_3839_3808_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_3807_3776_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_3775_3744_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_3743_3712_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_3711_3680_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_3679_3648_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_3647_3616_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_3615_3584_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_3583_3552_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_3551_3520_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_3519_3488_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_3487_3456_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_3455_3424_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_3423_3392_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_3391_3360_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_3359_3328_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_3327_3296_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_3295_3264_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_3263_3232_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_3231_3200_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_3199_3168_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_3167_3136_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_3135_3104_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_3103_3072_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_3071_3040_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_3039_3008_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_3007_2976_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_2975_2944_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_2943_2912_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_2911_2880_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_2879_2848_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_2847_2816_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_2815_2784_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_2783_2752_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_2751_2720_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_2719_2688_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_2687_2656_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_2655_2624_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_2623_2592_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_2591_2560_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_2559_2528_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_2527_2496_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_2495_2464_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_2463_2432_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_2431_2400_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_2399_2368_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_2367_2336_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_2335_2304_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_2303_2272_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_2271_2240_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_2239_2208_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_2207_2176_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_2175_2144_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_2143_2112_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_2111_2080_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_2079_2048_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_2047_2016_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_2015_1984_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_1983_1952_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_1951_1920_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_1919_1888_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_1887_1856_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_1855_1824_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_1823_1792_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_1791_1760_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_1759_1728_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_1727_1696_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_1695_1664_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_1663_1632_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_1631_1600_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_1599_1568_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_1567_1536_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_1535_1504_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_1503_1472_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_1471_1440_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_1439_1408_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_1407_1376_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_1375_1344_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_1343_1312_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_1311_1280_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_1279_1248_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_1247_1216_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_1215_1184_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_1183_1152_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_1151_1120_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_1119_1088_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_1087_1056_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_1055_1024_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_1023_992_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_991_960_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_959_928_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_927_896_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_895_864_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_863_832_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_831_800_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_799_768_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_767_736_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_735_704_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_703_672_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_671_640_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_639_608_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_607_576_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_575_544_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_543_512_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_511_480_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_479_448_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_447_416_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_415_384_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_383_352_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_351_320_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_319_288_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_287_256_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_255_224_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_223_192_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_191_160_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_159_128_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_127_96_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_95_64_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_63_32_lpi_2_dfm;
  reg [31:0] for_io_read_output_rsc_sdt_31_0_lpi_2_dfm;
  reg [31:0] for_mux_itm;
  wire [31:0] for_for_mul_1_cmx_sva_1;
  wire signed [36:0] nl_for_for_mul_1_cmx_sva_1;
  wire reg_output_rsc_1_31_output_or_cse;

  wire[0:0] and_660_nl;
  wire[0:0] and_666_nl;
  wire[0:0] and_672_nl;
  wire[0:0] and_678_nl;
  wire[0:0] and_684_nl;
  wire[0:0] and_690_nl;
  wire[0:0] and_696_nl;
  wire[0:0] and_702_nl;
  wire[0:0] and_708_nl;
  wire[0:0] and_714_nl;
  wire[0:0] and_720_nl;
  wire[0:0] and_726_nl;
  wire[0:0] and_732_nl;
  wire[0:0] and_738_nl;
  wire[0:0] and_744_nl;
  wire[0:0] and_750_nl;
  wire[0:0] and_756_nl;
  wire[0:0] and_762_nl;
  wire[0:0] and_768_nl;
  wire[0:0] and_774_nl;
  wire[0:0] and_780_nl;
  wire[0:0] and_786_nl;
  wire[0:0] and_792_nl;
  wire[0:0] and_798_nl;
  wire[0:0] and_804_nl;
  wire[0:0] and_810_nl;
  wire[0:0] and_816_nl;
  wire[0:0] and_822_nl;
  wire[0:0] and_828_nl;
  wire[0:0] and_834_nl;
  wire[0:0] and_840_nl;
  wire[0:0] and_846_nl;
  wire[0:0] and_852_nl;
  wire[0:0] and_858_nl;
  wire[0:0] and_864_nl;
  wire[0:0] and_870_nl;
  wire[0:0] and_876_nl;
  wire[0:0] and_882_nl;
  wire[0:0] and_888_nl;
  wire[0:0] and_894_nl;
  wire[0:0] and_900_nl;
  wire[0:0] and_906_nl;
  wire[0:0] and_912_nl;
  wire[0:0] and_918_nl;
  wire[0:0] and_924_nl;
  wire[0:0] and_930_nl;
  wire[0:0] and_936_nl;
  wire[0:0] and_942_nl;
  wire[0:0] and_948_nl;
  wire[0:0] and_954_nl;
  wire[0:0] and_960_nl;
  wire[0:0] and_966_nl;
  wire[0:0] and_972_nl;
  wire[0:0] and_978_nl;
  wire[0:0] and_984_nl;
  wire[0:0] and_990_nl;
  wire[0:0] and_996_nl;
  wire[0:0] and_1002_nl;
  wire[0:0] and_1008_nl;
  wire[0:0] and_1014_nl;
  wire[0:0] and_1020_nl;
  wire[0:0] and_1026_nl;
  wire[0:0] and_1032_nl;
  wire[0:0] and_1038_nl;
  wire[0:0] and_1044_nl;
  wire[0:0] and_1050_nl;
  wire[0:0] and_1056_nl;
  wire[0:0] and_1062_nl;
  wire[0:0] and_1068_nl;
  wire[0:0] and_1074_nl;
  wire[0:0] and_1080_nl;
  wire[0:0] and_1086_nl;
  wire[0:0] and_1092_nl;
  wire[0:0] and_1098_nl;
  wire[0:0] and_1104_nl;
  wire[0:0] and_1110_nl;
  wire[0:0] and_1116_nl;
  wire[0:0] and_1122_nl;
  wire[0:0] and_1128_nl;
  wire[0:0] and_1134_nl;
  wire[0:0] and_1140_nl;
  wire[0:0] and_1146_nl;
  wire[0:0] and_1152_nl;
  wire[0:0] and_1158_nl;
  wire[0:0] and_1164_nl;
  wire[0:0] and_1170_nl;
  wire[0:0] and_1176_nl;
  wire[0:0] and_1182_nl;
  wire[0:0] and_1188_nl;
  wire[0:0] and_1194_nl;
  wire[0:0] and_1200_nl;
  wire[0:0] and_1206_nl;
  wire[0:0] and_1212_nl;
  wire[0:0] and_1218_nl;
  wire[0:0] and_1224_nl;
  wire[0:0] and_1230_nl;
  wire[0:0] and_1236_nl;
  wire[0:0] and_1242_nl;
  wire[0:0] and_1248_nl;
  wire[0:0] and_1254_nl;
  wire[0:0] and_1260_nl;
  wire[0:0] and_1266_nl;
  wire[0:0] and_1272_nl;
  wire[0:0] and_1278_nl;
  wire[0:0] and_1284_nl;
  wire[0:0] and_1290_nl;
  wire[0:0] and_1296_nl;
  wire[0:0] and_1302_nl;
  wire[0:0] and_1308_nl;
  wire[0:0] and_1314_nl;
  wire[0:0] and_1320_nl;
  wire[0:0] and_1326_nl;
  wire[0:0] and_1332_nl;
  wire[0:0] and_1338_nl;
  wire[0:0] and_1344_nl;
  wire[0:0] and_1350_nl;
  wire[0:0] and_1356_nl;
  wire[0:0] and_1362_nl;
  wire[0:0] and_1368_nl;
  wire[0:0] and_1374_nl;
  wire[0:0] and_1380_nl;
  wire[0:0] and_1386_nl;
  wire[0:0] and_1392_nl;
  wire[0:0] and_1398_nl;
  wire[0:0] and_1404_nl;
  wire[0:0] and_1410_nl;
  wire[0:0] and_1416_nl;
  wire[0:0] for_and_253_nl;
  wire[0:0] for_and_251_nl;
  wire[0:0] for_and_249_nl;
  wire[0:0] for_and_247_nl;
  wire[0:0] for_and_245_nl;
  wire[0:0] for_and_243_nl;
  wire[0:0] for_and_241_nl;
  wire[0:0] for_and_239_nl;
  wire[0:0] for_and_237_nl;
  wire[0:0] for_and_235_nl;
  wire[0:0] for_and_233_nl;
  wire[0:0] for_and_231_nl;
  wire[0:0] for_and_229_nl;
  wire[0:0] for_and_227_nl;
  wire[0:0] for_and_225_nl;
  wire[0:0] for_and_223_nl;
  wire[0:0] for_and_221_nl;
  wire[0:0] for_and_219_nl;
  wire[0:0] for_and_217_nl;
  wire[0:0] for_and_215_nl;
  wire[0:0] for_and_213_nl;
  wire[0:0] for_and_211_nl;
  wire[0:0] for_and_209_nl;
  wire[0:0] for_and_207_nl;
  wire[0:0] for_and_205_nl;
  wire[0:0] for_and_203_nl;
  wire[0:0] for_and_201_nl;
  wire[0:0] for_and_199_nl;
  wire[0:0] for_and_197_nl;
  wire[0:0] for_and_195_nl;
  wire[0:0] for_and_193_nl;
  wire[0:0] for_and_191_nl;
  wire[0:0] for_and_189_nl;
  wire[0:0] for_and_187_nl;
  wire[0:0] for_and_185_nl;
  wire[0:0] for_and_183_nl;
  wire[0:0] for_and_181_nl;
  wire[0:0] for_and_179_nl;
  wire[0:0] for_and_177_nl;
  wire[0:0] for_and_175_nl;
  wire[0:0] for_and_173_nl;
  wire[0:0] for_and_171_nl;
  wire[0:0] for_and_169_nl;
  wire[0:0] for_and_167_nl;
  wire[0:0] for_and_165_nl;
  wire[0:0] for_and_163_nl;
  wire[0:0] for_and_161_nl;
  wire[0:0] for_and_159_nl;
  wire[0:0] for_and_157_nl;
  wire[0:0] for_and_155_nl;
  wire[0:0] for_and_153_nl;
  wire[0:0] for_and_151_nl;
  wire[0:0] for_and_149_nl;
  wire[0:0] for_and_147_nl;
  wire[0:0] for_and_145_nl;
  wire[0:0] for_and_143_nl;
  wire[0:0] for_and_141_nl;
  wire[0:0] for_and_139_nl;
  wire[0:0] for_and_137_nl;
  wire[0:0] for_and_135_nl;
  wire[0:0] for_and_133_nl;
  wire[0:0] for_and_131_nl;
  wire[0:0] for_and_129_nl;
  wire[0:0] for_and_127_nl;
  wire[0:0] for_and_125_nl;
  wire[0:0] for_and_123_nl;
  wire[0:0] for_and_121_nl;
  wire[0:0] for_and_119_nl;
  wire[0:0] for_and_117_nl;
  wire[0:0] for_and_115_nl;
  wire[0:0] for_and_113_nl;
  wire[0:0] for_and_111_nl;
  wire[0:0] for_and_109_nl;
  wire[0:0] for_and_107_nl;
  wire[0:0] for_and_105_nl;
  wire[0:0] for_and_103_nl;
  wire[0:0] for_and_101_nl;
  wire[0:0] for_and_99_nl;
  wire[0:0] for_and_97_nl;
  wire[0:0] for_and_95_nl;
  wire[0:0] for_and_93_nl;
  wire[0:0] for_and_91_nl;
  wire[0:0] for_and_89_nl;
  wire[0:0] for_and_87_nl;
  wire[0:0] for_and_85_nl;
  wire[0:0] for_and_83_nl;
  wire[0:0] for_and_81_nl;
  wire[0:0] for_and_79_nl;
  wire[0:0] for_and_77_nl;
  wire[0:0] for_and_75_nl;
  wire[0:0] for_and_73_nl;
  wire[0:0] for_and_71_nl;
  wire[0:0] for_and_69_nl;
  wire[0:0] for_and_67_nl;
  wire[0:0] for_and_65_nl;
  wire[0:0] for_and_63_nl;
  wire[0:0] for_and_61_nl;
  wire[0:0] for_and_59_nl;
  wire[0:0] for_and_57_nl;
  wire[0:0] for_and_55_nl;
  wire[0:0] for_and_53_nl;
  wire[0:0] for_and_51_nl;
  wire[0:0] for_and_49_nl;
  wire[0:0] for_and_47_nl;
  wire[0:0] for_and_45_nl;
  wire[0:0] for_and_43_nl;
  wire[0:0] for_and_41_nl;
  wire[0:0] for_and_39_nl;
  wire[0:0] for_and_37_nl;
  wire[0:0] for_and_35_nl;
  wire[0:0] for_and_33_nl;
  wire[0:0] for_and_31_nl;
  wire[0:0] for_and_29_nl;
  wire[0:0] for_and_27_nl;
  wire[0:0] for_and_25_nl;
  wire[0:0] for_and_23_nl;
  wire[0:0] for_and_21_nl;
  wire[0:0] for_and_19_nl;
  wire[0:0] for_and_17_nl;
  wire[0:0] for_and_15_nl;
  wire[0:0] for_and_13_nl;
  wire[0:0] for_and_11_nl;
  wire[0:0] for_and_9_nl;
  wire[0:0] for_and_7_nl;
  wire[0:0] for_and_5_nl;
  wire[0:0] for_and_3_nl;
  wire[0:0] for_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [4095:0] nl_output_rsci_idat;
  assign nl_output_rsci_idat = {output_rsci_idat_4095_4064 , output_rsci_idat_4063_4032
      , output_rsci_idat_4031_4000 , output_rsci_idat_3999_3968 , output_rsci_idat_3967_3936
      , output_rsci_idat_3935_3904 , output_rsci_idat_3903_3872 , output_rsci_idat_3871_3840
      , output_rsci_idat_3839_3808 , output_rsci_idat_3807_3776 , output_rsci_idat_3775_3744
      , output_rsci_idat_3743_3712 , output_rsci_idat_3711_3680 , output_rsci_idat_3679_3648
      , output_rsci_idat_3647_3616 , output_rsci_idat_3615_3584 , output_rsci_idat_3583_3552
      , output_rsci_idat_3551_3520 , output_rsci_idat_3519_3488 , output_rsci_idat_3487_3456
      , output_rsci_idat_3455_3424 , output_rsci_idat_3423_3392 , output_rsci_idat_3391_3360
      , output_rsci_idat_3359_3328 , output_rsci_idat_3327_3296 , output_rsci_idat_3295_3264
      , output_rsci_idat_3263_3232 , output_rsci_idat_3231_3200 , output_rsci_idat_3199_3168
      , output_rsci_idat_3167_3136 , output_rsci_idat_3135_3104 , output_rsci_idat_3103_3072
      , output_rsci_idat_3071_3040 , output_rsci_idat_3039_3008 , output_rsci_idat_3007_2976
      , output_rsci_idat_2975_2944 , output_rsci_idat_2943_2912 , output_rsci_idat_2911_2880
      , output_rsci_idat_2879_2848 , output_rsci_idat_2847_2816 , output_rsci_idat_2815_2784
      , output_rsci_idat_2783_2752 , output_rsci_idat_2751_2720 , output_rsci_idat_2719_2688
      , output_rsci_idat_2687_2656 , output_rsci_idat_2655_2624 , output_rsci_idat_2623_2592
      , output_rsci_idat_2591_2560 , output_rsci_idat_2559_2528 , output_rsci_idat_2527_2496
      , output_rsci_idat_2495_2464 , output_rsci_idat_2463_2432 , output_rsci_idat_2431_2400
      , output_rsci_idat_2399_2368 , output_rsci_idat_2367_2336 , output_rsci_idat_2335_2304
      , output_rsci_idat_2303_2272 , output_rsci_idat_2271_2240 , output_rsci_idat_2239_2208
      , output_rsci_idat_2207_2176 , output_rsci_idat_2175_2144 , output_rsci_idat_2143_2112
      , output_rsci_idat_2111_2080 , output_rsci_idat_2079_2048 , output_rsci_idat_2047_2016
      , output_rsci_idat_2015_1984 , output_rsci_idat_1983_1952 , output_rsci_idat_1951_1920
      , output_rsci_idat_1919_1888 , output_rsci_idat_1887_1856 , output_rsci_idat_1855_1824
      , output_rsci_idat_1823_1792 , output_rsci_idat_1791_1760 , output_rsci_idat_1759_1728
      , output_rsci_idat_1727_1696 , output_rsci_idat_1695_1664 , output_rsci_idat_1663_1632
      , output_rsci_idat_1631_1600 , output_rsci_idat_1599_1568 , output_rsci_idat_1567_1536
      , output_rsci_idat_1535_1504 , output_rsci_idat_1503_1472 , output_rsci_idat_1471_1440
      , output_rsci_idat_1439_1408 , output_rsci_idat_1407_1376 , output_rsci_idat_1375_1344
      , output_rsci_idat_1343_1312 , output_rsci_idat_1311_1280 , output_rsci_idat_1279_1248
      , output_rsci_idat_1247_1216 , output_rsci_idat_1215_1184 , output_rsci_idat_1183_1152
      , output_rsci_idat_1151_1120 , output_rsci_idat_1119_1088 , output_rsci_idat_1087_1056
      , output_rsci_idat_1055_1024 , output_rsci_idat_1023_992 , output_rsci_idat_991_960
      , output_rsci_idat_959_928 , output_rsci_idat_927_896 , output_rsci_idat_895_864
      , output_rsci_idat_863_832 , output_rsci_idat_831_800 , output_rsci_idat_799_768
      , output_rsci_idat_767_736 , output_rsci_idat_735_704 , output_rsci_idat_703_672
      , output_rsci_idat_671_640 , output_rsci_idat_639_608 , output_rsci_idat_607_576
      , output_rsci_idat_575_544 , output_rsci_idat_543_512 , output_rsci_idat_511_480
      , output_rsci_idat_479_448 , output_rsci_idat_447_416 , output_rsci_idat_415_384
      , output_rsci_idat_383_352 , output_rsci_idat_351_320 , output_rsci_idat_319_288
      , output_rsci_idat_287_256 , output_rsci_idat_255_224 , output_rsci_idat_223_192
      , output_rsci_idat_191_160 , output_rsci_idat_159_128 , output_rsci_idat_127_96
      , output_rsci_idat_95_64 , output_rsci_idat_63_32 , output_rsci_idat_31_0};
  wire [0:0] nl_fir_core_core_fsm_inst_for_C_2_tr0;
  assign nl_fir_core_core_fsm_inst_for_C_2_tr0 = i_7_0_sva_1[7];
  ccs_in_v1 #(.rscid(32'sd1),
  .width(32'sd4096)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  ccs_out_v1 #(.rscid(32'sd2),
  .width(32'sd4096)) output_rsci (
      .idat(nl_output_rsci_idat[4095:0]),
      .dat(output_rsc_dat)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) input_rsc_triosy_obj (
      .ld(reg_output_rsc_triosy_obj_ld_cse),
      .lz(input_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) output_rsc_triosy_obj (
      .ld(reg_output_rsc_triosy_obj_ld_cse),
      .lz(output_rsc_triosy_lz)
    );
  fir_core_core_fsm fir_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output),
      .for_C_2_tr0(nl_fir_core_core_fsm_inst_for_C_2_tr0[0:0])
    );
  assign reg_output_rsc_1_31_output_or_cse = (fsm_output[3]) | (fsm_output[0]);
  assign output_output_mux_cse = MUX_v_32_2_2(output_rsc_1_31_0_lpi_2, for_for_mul_1_cmx_sva_1,
      or_tmp_259);
  assign nl_for_for_mul_1_cmx_sva_1 = $signed(for_mux_itm) * $signed(5'b01101);
  assign for_for_mul_1_cmx_sva_1 = nl_for_for_mul_1_cmx_sva_1[31:0];
  assign for_or_tmp = ((i_7_0_sva_6_0[0]) & for_nor_itm) | ((i_7_0_sva_6_0[1]) &
      for_nor_1_itm) | for_equal_tmp_3 | ((i_7_0_sva_6_0[2]) & for_nor_3_itm) | for_equal_tmp_5
      | for_equal_tmp_6 | for_equal_tmp_7 | ((i_7_0_sva_6_0[3]) & for_nor_7_itm)
      | for_equal_tmp_9 | for_equal_tmp_10 | for_equal_tmp_11 | for_equal_tmp_12
      | for_equal_tmp_13 | for_equal_tmp_14 | for_equal_tmp_15 | ((i_7_0_sva_6_0[4])
      & for_nor_15_itm) | for_equal_tmp_17 | for_equal_tmp_18 | for_equal_tmp_19
      | for_equal_tmp_20 | for_equal_tmp_21 | for_equal_tmp_22 | for_equal_tmp_23
      | for_equal_tmp_24 | for_equal_tmp_25 | for_equal_tmp_26 | for_equal_tmp_27
      | for_equal_tmp_28 | for_equal_tmp_29 | for_equal_tmp_30 | for_equal_tmp_31
      | ((i_7_0_sva_6_0[5]) & for_nor_31_itm) | for_equal_tmp_33 | for_equal_tmp_34
      | for_equal_tmp_35 | for_equal_tmp_36 | for_equal_tmp_37 | for_equal_tmp_38
      | for_equal_tmp_39 | for_equal_tmp_40 | for_equal_tmp_41 | for_equal_tmp_42
      | for_equal_tmp_43 | for_equal_tmp_44 | for_equal_tmp_45 | for_equal_tmp_46
      | for_equal_tmp_47 | for_equal_tmp_48 | for_equal_tmp_49 | for_equal_tmp_50
      | for_equal_tmp_51 | for_equal_tmp_52 | for_equal_tmp_53 | for_equal_tmp_54
      | for_equal_tmp_55 | for_equal_tmp_56 | for_equal_tmp_57 | for_equal_tmp_58
      | for_equal_tmp_59 | for_equal_tmp_60 | for_equal_tmp_61 | for_equal_tmp_62
      | for_equal_tmp_63 | ((i_7_0_sva_6_0[6]) & for_nor_62_itm) | for_equal_tmp_65
      | for_equal_tmp_66 | for_equal_tmp_67 | for_equal_tmp_68 | for_equal_tmp_69
      | for_equal_tmp_70 | for_equal_tmp_71 | for_equal_tmp_72 | for_equal_tmp_73
      | for_equal_tmp_74 | for_equal_tmp_75 | for_equal_tmp_76 | for_equal_tmp_77
      | for_equal_tmp_78 | for_equal_tmp_79 | for_equal_tmp_80 | for_equal_tmp_81
      | for_equal_tmp_82 | for_equal_tmp_83 | for_equal_tmp_84 | for_equal_tmp_85
      | for_equal_tmp_86 | for_equal_tmp_87 | for_equal_tmp_88 | for_equal_tmp_89
      | for_equal_tmp_90 | for_equal_tmp_91 | for_equal_tmp_92 | for_equal_tmp_93
      | for_equal_tmp_94 | for_equal_tmp_95 | for_equal_tmp_96 | for_equal_tmp_97
      | for_equal_tmp_98 | for_equal_tmp_99 | for_equal_tmp_100 | for_equal_tmp_101
      | for_equal_tmp_102 | for_equal_tmp_103 | for_equal_tmp_104 | for_equal_tmp_105
      | for_equal_tmp_106 | for_equal_tmp_107 | for_equal_tmp_108 | for_equal_tmp_109
      | for_equal_tmp_110 | for_equal_tmp_111 | for_equal_tmp_112 | for_equal_tmp_113
      | for_equal_tmp_114 | for_equal_tmp_115 | for_equal_tmp_116 | for_equal_tmp_117
      | for_equal_tmp_118 | for_equal_tmp_119 | for_equal_tmp_120 | for_equal_tmp_121
      | for_equal_tmp_122 | for_equal_tmp_123 | for_equal_tmp_124 | for_equal_tmp_125
      | for_equal_tmp_126 | for_equal_tmp_127;
  assign or_dcpl_330 = ~((i_7_0_sva_6_0[0]) & for_nor_itm);
  assign or_dcpl_331 = ~((i_7_0_sva_6_0[1]) & for_nor_1_itm);
  assign or_dcpl_332 = ~((i_7_0_sva_6_0[2]) & for_nor_3_itm);
  assign or_dcpl_333 = ~((i_7_0_sva_6_0[3]) & for_nor_7_itm);
  assign or_dcpl_334 = ~((i_7_0_sva_6_0[4]) & for_nor_15_itm);
  assign or_dcpl_335 = ~((i_7_0_sva_6_0[5]) & for_nor_31_itm);
  assign or_dcpl_336 = ~(for_nor_62_itm & (i_7_0_sva_6_0[6]));
  assign or_tmp_259 = (~ for_or_tmp) & (fsm_output[2]);
  assign or_tmp_643 = (fsm_output[4:3]!=2'b00);
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsc_1_31_0_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_63_32_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_95_64_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_127_96_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_159_128_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_191_160_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_223_192_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_255_224_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_287_256_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_319_288_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_351_320_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_383_352_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_415_384_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_447_416_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_479_448_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_511_480_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_543_512_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_575_544_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_607_576_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_639_608_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_671_640_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_703_672_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_735_704_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_767_736_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_799_768_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_831_800_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_863_832_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_895_864_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_927_896_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_959_928_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_991_960_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_1023_992_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_1055_1024_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_1087_1056_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_1119_1088_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_1151_1120_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_1183_1152_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_1215_1184_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_1247_1216_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_1279_1248_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_1311_1280_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_1343_1312_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_1375_1344_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_1407_1376_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_1439_1408_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_1471_1440_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_1503_1472_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_1535_1504_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_1567_1536_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_1599_1568_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_1631_1600_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_1663_1632_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_1695_1664_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_1727_1696_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_1759_1728_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_1791_1760_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_1823_1792_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_1855_1824_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_1887_1856_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_1919_1888_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_1951_1920_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_1983_1952_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_2015_1984_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_2047_2016_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_2079_2048_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_2111_2080_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_2143_2112_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_2175_2144_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_2207_2176_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_2239_2208_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_2271_2240_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_2303_2272_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_2335_2304_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_2367_2336_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_2399_2368_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_2431_2400_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_2463_2432_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_2495_2464_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_2527_2496_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_2559_2528_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_2591_2560_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_2623_2592_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_2655_2624_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_2687_2656_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_2719_2688_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_2751_2720_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_2783_2752_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_2815_2784_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_2847_2816_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_2879_2848_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_2911_2880_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_2943_2912_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_2975_2944_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_3007_2976_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_3039_3008_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_3071_3040_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_3103_3072_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_3135_3104_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_3167_3136_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_3199_3168_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_3231_3200_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_3263_3232_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_3295_3264_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_3327_3296_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_3359_3328_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_3391_3360_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_3423_3392_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_3455_3424_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_3487_3456_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_3519_3488_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_3551_3520_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_3583_3552_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_3615_3584_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_3647_3616_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_3679_3648_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_3711_3680_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_3743_3712_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_3775_3744_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_3807_3776_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_3839_3808_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_3871_3840_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_3903_3872_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_3935_3904_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_3967_3936_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_3999_3968_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_4031_4000_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_4063_4032_lpi_2 <= 32'b00000000000000000000000000000000;
      output_rsc_1_4095_4064_lpi_2 <= 32'b00000000000000000000000000000000;
      i_7_0_sva_6_0 <= 7'b0000000;
    end
    else if ( reg_output_rsc_1_31_output_or_cse ) begin
      output_rsc_1_31_0_lpi_2 <= for_io_read_output_rsc_sdt_31_0_lpi_2_dfm;
      output_rsc_1_63_32_lpi_2 <= for_io_read_output_rsc_sdt_63_32_lpi_2_dfm;
      output_rsc_1_95_64_lpi_2 <= for_io_read_output_rsc_sdt_95_64_lpi_2_dfm;
      output_rsc_1_127_96_lpi_2 <= for_io_read_output_rsc_sdt_127_96_lpi_2_dfm;
      output_rsc_1_159_128_lpi_2 <= for_io_read_output_rsc_sdt_159_128_lpi_2_dfm;
      output_rsc_1_191_160_lpi_2 <= for_io_read_output_rsc_sdt_191_160_lpi_2_dfm;
      output_rsc_1_223_192_lpi_2 <= for_io_read_output_rsc_sdt_223_192_lpi_2_dfm;
      output_rsc_1_255_224_lpi_2 <= for_io_read_output_rsc_sdt_255_224_lpi_2_dfm;
      output_rsc_1_287_256_lpi_2 <= for_io_read_output_rsc_sdt_287_256_lpi_2_dfm;
      output_rsc_1_319_288_lpi_2 <= for_io_read_output_rsc_sdt_319_288_lpi_2_dfm;
      output_rsc_1_351_320_lpi_2 <= for_io_read_output_rsc_sdt_351_320_lpi_2_dfm;
      output_rsc_1_383_352_lpi_2 <= for_io_read_output_rsc_sdt_383_352_lpi_2_dfm;
      output_rsc_1_415_384_lpi_2 <= for_io_read_output_rsc_sdt_415_384_lpi_2_dfm;
      output_rsc_1_447_416_lpi_2 <= for_io_read_output_rsc_sdt_447_416_lpi_2_dfm;
      output_rsc_1_479_448_lpi_2 <= for_io_read_output_rsc_sdt_479_448_lpi_2_dfm;
      output_rsc_1_511_480_lpi_2 <= for_io_read_output_rsc_sdt_511_480_lpi_2_dfm;
      output_rsc_1_543_512_lpi_2 <= for_io_read_output_rsc_sdt_543_512_lpi_2_dfm;
      output_rsc_1_575_544_lpi_2 <= for_io_read_output_rsc_sdt_575_544_lpi_2_dfm;
      output_rsc_1_607_576_lpi_2 <= for_io_read_output_rsc_sdt_607_576_lpi_2_dfm;
      output_rsc_1_639_608_lpi_2 <= for_io_read_output_rsc_sdt_639_608_lpi_2_dfm;
      output_rsc_1_671_640_lpi_2 <= for_io_read_output_rsc_sdt_671_640_lpi_2_dfm;
      output_rsc_1_703_672_lpi_2 <= for_io_read_output_rsc_sdt_703_672_lpi_2_dfm;
      output_rsc_1_735_704_lpi_2 <= for_io_read_output_rsc_sdt_735_704_lpi_2_dfm;
      output_rsc_1_767_736_lpi_2 <= for_io_read_output_rsc_sdt_767_736_lpi_2_dfm;
      output_rsc_1_799_768_lpi_2 <= for_io_read_output_rsc_sdt_799_768_lpi_2_dfm;
      output_rsc_1_831_800_lpi_2 <= for_io_read_output_rsc_sdt_831_800_lpi_2_dfm;
      output_rsc_1_863_832_lpi_2 <= for_io_read_output_rsc_sdt_863_832_lpi_2_dfm;
      output_rsc_1_895_864_lpi_2 <= for_io_read_output_rsc_sdt_895_864_lpi_2_dfm;
      output_rsc_1_927_896_lpi_2 <= for_io_read_output_rsc_sdt_927_896_lpi_2_dfm;
      output_rsc_1_959_928_lpi_2 <= for_io_read_output_rsc_sdt_959_928_lpi_2_dfm;
      output_rsc_1_991_960_lpi_2 <= for_io_read_output_rsc_sdt_991_960_lpi_2_dfm;
      output_rsc_1_1023_992_lpi_2 <= for_io_read_output_rsc_sdt_1023_992_lpi_2_dfm;
      output_rsc_1_1055_1024_lpi_2 <= for_io_read_output_rsc_sdt_1055_1024_lpi_2_dfm;
      output_rsc_1_1087_1056_lpi_2 <= for_io_read_output_rsc_sdt_1087_1056_lpi_2_dfm;
      output_rsc_1_1119_1088_lpi_2 <= for_io_read_output_rsc_sdt_1119_1088_lpi_2_dfm;
      output_rsc_1_1151_1120_lpi_2 <= for_io_read_output_rsc_sdt_1151_1120_lpi_2_dfm;
      output_rsc_1_1183_1152_lpi_2 <= for_io_read_output_rsc_sdt_1183_1152_lpi_2_dfm;
      output_rsc_1_1215_1184_lpi_2 <= for_io_read_output_rsc_sdt_1215_1184_lpi_2_dfm;
      output_rsc_1_1247_1216_lpi_2 <= for_io_read_output_rsc_sdt_1247_1216_lpi_2_dfm;
      output_rsc_1_1279_1248_lpi_2 <= for_io_read_output_rsc_sdt_1279_1248_lpi_2_dfm;
      output_rsc_1_1311_1280_lpi_2 <= for_io_read_output_rsc_sdt_1311_1280_lpi_2_dfm;
      output_rsc_1_1343_1312_lpi_2 <= for_io_read_output_rsc_sdt_1343_1312_lpi_2_dfm;
      output_rsc_1_1375_1344_lpi_2 <= for_io_read_output_rsc_sdt_1375_1344_lpi_2_dfm;
      output_rsc_1_1407_1376_lpi_2 <= for_io_read_output_rsc_sdt_1407_1376_lpi_2_dfm;
      output_rsc_1_1439_1408_lpi_2 <= for_io_read_output_rsc_sdt_1439_1408_lpi_2_dfm;
      output_rsc_1_1471_1440_lpi_2 <= for_io_read_output_rsc_sdt_1471_1440_lpi_2_dfm;
      output_rsc_1_1503_1472_lpi_2 <= for_io_read_output_rsc_sdt_1503_1472_lpi_2_dfm;
      output_rsc_1_1535_1504_lpi_2 <= for_io_read_output_rsc_sdt_1535_1504_lpi_2_dfm;
      output_rsc_1_1567_1536_lpi_2 <= for_io_read_output_rsc_sdt_1567_1536_lpi_2_dfm;
      output_rsc_1_1599_1568_lpi_2 <= for_io_read_output_rsc_sdt_1599_1568_lpi_2_dfm;
      output_rsc_1_1631_1600_lpi_2 <= for_io_read_output_rsc_sdt_1631_1600_lpi_2_dfm;
      output_rsc_1_1663_1632_lpi_2 <= for_io_read_output_rsc_sdt_1663_1632_lpi_2_dfm;
      output_rsc_1_1695_1664_lpi_2 <= for_io_read_output_rsc_sdt_1695_1664_lpi_2_dfm;
      output_rsc_1_1727_1696_lpi_2 <= for_io_read_output_rsc_sdt_1727_1696_lpi_2_dfm;
      output_rsc_1_1759_1728_lpi_2 <= for_io_read_output_rsc_sdt_1759_1728_lpi_2_dfm;
      output_rsc_1_1791_1760_lpi_2 <= for_io_read_output_rsc_sdt_1791_1760_lpi_2_dfm;
      output_rsc_1_1823_1792_lpi_2 <= for_io_read_output_rsc_sdt_1823_1792_lpi_2_dfm;
      output_rsc_1_1855_1824_lpi_2 <= for_io_read_output_rsc_sdt_1855_1824_lpi_2_dfm;
      output_rsc_1_1887_1856_lpi_2 <= for_io_read_output_rsc_sdt_1887_1856_lpi_2_dfm;
      output_rsc_1_1919_1888_lpi_2 <= for_io_read_output_rsc_sdt_1919_1888_lpi_2_dfm;
      output_rsc_1_1951_1920_lpi_2 <= for_io_read_output_rsc_sdt_1951_1920_lpi_2_dfm;
      output_rsc_1_1983_1952_lpi_2 <= for_io_read_output_rsc_sdt_1983_1952_lpi_2_dfm;
      output_rsc_1_2015_1984_lpi_2 <= for_io_read_output_rsc_sdt_2015_1984_lpi_2_dfm;
      output_rsc_1_2047_2016_lpi_2 <= for_io_read_output_rsc_sdt_2047_2016_lpi_2_dfm;
      output_rsc_1_2079_2048_lpi_2 <= for_io_read_output_rsc_sdt_2079_2048_lpi_2_dfm;
      output_rsc_1_2111_2080_lpi_2 <= for_io_read_output_rsc_sdt_2111_2080_lpi_2_dfm;
      output_rsc_1_2143_2112_lpi_2 <= for_io_read_output_rsc_sdt_2143_2112_lpi_2_dfm;
      output_rsc_1_2175_2144_lpi_2 <= for_io_read_output_rsc_sdt_2175_2144_lpi_2_dfm;
      output_rsc_1_2207_2176_lpi_2 <= for_io_read_output_rsc_sdt_2207_2176_lpi_2_dfm;
      output_rsc_1_2239_2208_lpi_2 <= for_io_read_output_rsc_sdt_2239_2208_lpi_2_dfm;
      output_rsc_1_2271_2240_lpi_2 <= for_io_read_output_rsc_sdt_2271_2240_lpi_2_dfm;
      output_rsc_1_2303_2272_lpi_2 <= for_io_read_output_rsc_sdt_2303_2272_lpi_2_dfm;
      output_rsc_1_2335_2304_lpi_2 <= for_io_read_output_rsc_sdt_2335_2304_lpi_2_dfm;
      output_rsc_1_2367_2336_lpi_2 <= for_io_read_output_rsc_sdt_2367_2336_lpi_2_dfm;
      output_rsc_1_2399_2368_lpi_2 <= for_io_read_output_rsc_sdt_2399_2368_lpi_2_dfm;
      output_rsc_1_2431_2400_lpi_2 <= for_io_read_output_rsc_sdt_2431_2400_lpi_2_dfm;
      output_rsc_1_2463_2432_lpi_2 <= for_io_read_output_rsc_sdt_2463_2432_lpi_2_dfm;
      output_rsc_1_2495_2464_lpi_2 <= for_io_read_output_rsc_sdt_2495_2464_lpi_2_dfm;
      output_rsc_1_2527_2496_lpi_2 <= for_io_read_output_rsc_sdt_2527_2496_lpi_2_dfm;
      output_rsc_1_2559_2528_lpi_2 <= for_io_read_output_rsc_sdt_2559_2528_lpi_2_dfm;
      output_rsc_1_2591_2560_lpi_2 <= for_io_read_output_rsc_sdt_2591_2560_lpi_2_dfm;
      output_rsc_1_2623_2592_lpi_2 <= for_io_read_output_rsc_sdt_2623_2592_lpi_2_dfm;
      output_rsc_1_2655_2624_lpi_2 <= for_io_read_output_rsc_sdt_2655_2624_lpi_2_dfm;
      output_rsc_1_2687_2656_lpi_2 <= for_io_read_output_rsc_sdt_2687_2656_lpi_2_dfm;
      output_rsc_1_2719_2688_lpi_2 <= for_io_read_output_rsc_sdt_2719_2688_lpi_2_dfm;
      output_rsc_1_2751_2720_lpi_2 <= for_io_read_output_rsc_sdt_2751_2720_lpi_2_dfm;
      output_rsc_1_2783_2752_lpi_2 <= for_io_read_output_rsc_sdt_2783_2752_lpi_2_dfm;
      output_rsc_1_2815_2784_lpi_2 <= for_io_read_output_rsc_sdt_2815_2784_lpi_2_dfm;
      output_rsc_1_2847_2816_lpi_2 <= for_io_read_output_rsc_sdt_2847_2816_lpi_2_dfm;
      output_rsc_1_2879_2848_lpi_2 <= for_io_read_output_rsc_sdt_2879_2848_lpi_2_dfm;
      output_rsc_1_2911_2880_lpi_2 <= for_io_read_output_rsc_sdt_2911_2880_lpi_2_dfm;
      output_rsc_1_2943_2912_lpi_2 <= for_io_read_output_rsc_sdt_2943_2912_lpi_2_dfm;
      output_rsc_1_2975_2944_lpi_2 <= for_io_read_output_rsc_sdt_2975_2944_lpi_2_dfm;
      output_rsc_1_3007_2976_lpi_2 <= for_io_read_output_rsc_sdt_3007_2976_lpi_2_dfm;
      output_rsc_1_3039_3008_lpi_2 <= for_io_read_output_rsc_sdt_3039_3008_lpi_2_dfm;
      output_rsc_1_3071_3040_lpi_2 <= for_io_read_output_rsc_sdt_3071_3040_lpi_2_dfm;
      output_rsc_1_3103_3072_lpi_2 <= for_io_read_output_rsc_sdt_3103_3072_lpi_2_dfm;
      output_rsc_1_3135_3104_lpi_2 <= for_io_read_output_rsc_sdt_3135_3104_lpi_2_dfm;
      output_rsc_1_3167_3136_lpi_2 <= for_io_read_output_rsc_sdt_3167_3136_lpi_2_dfm;
      output_rsc_1_3199_3168_lpi_2 <= for_io_read_output_rsc_sdt_3199_3168_lpi_2_dfm;
      output_rsc_1_3231_3200_lpi_2 <= for_io_read_output_rsc_sdt_3231_3200_lpi_2_dfm;
      output_rsc_1_3263_3232_lpi_2 <= for_io_read_output_rsc_sdt_3263_3232_lpi_2_dfm;
      output_rsc_1_3295_3264_lpi_2 <= for_io_read_output_rsc_sdt_3295_3264_lpi_2_dfm;
      output_rsc_1_3327_3296_lpi_2 <= for_io_read_output_rsc_sdt_3327_3296_lpi_2_dfm;
      output_rsc_1_3359_3328_lpi_2 <= for_io_read_output_rsc_sdt_3359_3328_lpi_2_dfm;
      output_rsc_1_3391_3360_lpi_2 <= for_io_read_output_rsc_sdt_3391_3360_lpi_2_dfm;
      output_rsc_1_3423_3392_lpi_2 <= for_io_read_output_rsc_sdt_3423_3392_lpi_2_dfm;
      output_rsc_1_3455_3424_lpi_2 <= for_io_read_output_rsc_sdt_3455_3424_lpi_2_dfm;
      output_rsc_1_3487_3456_lpi_2 <= for_io_read_output_rsc_sdt_3487_3456_lpi_2_dfm;
      output_rsc_1_3519_3488_lpi_2 <= for_io_read_output_rsc_sdt_3519_3488_lpi_2_dfm;
      output_rsc_1_3551_3520_lpi_2 <= for_io_read_output_rsc_sdt_3551_3520_lpi_2_dfm;
      output_rsc_1_3583_3552_lpi_2 <= for_io_read_output_rsc_sdt_3583_3552_lpi_2_dfm;
      output_rsc_1_3615_3584_lpi_2 <= for_io_read_output_rsc_sdt_3615_3584_lpi_2_dfm;
      output_rsc_1_3647_3616_lpi_2 <= for_io_read_output_rsc_sdt_3647_3616_lpi_2_dfm;
      output_rsc_1_3679_3648_lpi_2 <= for_io_read_output_rsc_sdt_3679_3648_lpi_2_dfm;
      output_rsc_1_3711_3680_lpi_2 <= for_io_read_output_rsc_sdt_3711_3680_lpi_2_dfm;
      output_rsc_1_3743_3712_lpi_2 <= for_io_read_output_rsc_sdt_3743_3712_lpi_2_dfm;
      output_rsc_1_3775_3744_lpi_2 <= for_io_read_output_rsc_sdt_3775_3744_lpi_2_dfm;
      output_rsc_1_3807_3776_lpi_2 <= for_io_read_output_rsc_sdt_3807_3776_lpi_2_dfm;
      output_rsc_1_3839_3808_lpi_2 <= for_io_read_output_rsc_sdt_3839_3808_lpi_2_dfm;
      output_rsc_1_3871_3840_lpi_2 <= for_io_read_output_rsc_sdt_3871_3840_lpi_2_dfm;
      output_rsc_1_3903_3872_lpi_2 <= for_io_read_output_rsc_sdt_3903_3872_lpi_2_dfm;
      output_rsc_1_3935_3904_lpi_2 <= for_io_read_output_rsc_sdt_3935_3904_lpi_2_dfm;
      output_rsc_1_3967_3936_lpi_2 <= for_io_read_output_rsc_sdt_3967_3936_lpi_2_dfm;
      output_rsc_1_3999_3968_lpi_2 <= for_io_read_output_rsc_sdt_3999_3968_lpi_2_dfm;
      output_rsc_1_4031_4000_lpi_2 <= for_io_read_output_rsc_sdt_4031_4000_lpi_2_dfm;
      output_rsc_1_4063_4032_lpi_2 <= for_io_read_output_rsc_sdt_4063_4032_lpi_2_dfm;
      output_rsc_1_4095_4064_lpi_2 <= for_io_read_output_rsc_sdt_4095_4064_lpi_2_dfm;
      i_7_0_sva_6_0 <= MUX_v_7_2_2(7'b0000000, (i_7_0_sva_1[6:0]), (fsm_output[3]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_31_0 <= 32'b00000000000000000000000000000000;
    end
    else if ( (for_or_tmp & (fsm_output[2])) | or_tmp_259 ) begin
      output_rsci_idat_31_0 <= output_output_mux_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_63_32 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_63_32 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_63_32_lpi_2,
          and_660_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_95_64 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_95_64 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_95_64_lpi_2,
          and_666_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_127_96 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_127_96 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_127_96_lpi_2,
          and_672_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_159_128 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_159_128 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_159_128_lpi_2,
          and_678_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_191_160 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_191_160 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_191_160_lpi_2,
          and_684_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_223_192 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_223_192 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_223_192_lpi_2,
          and_690_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_255_224 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_255_224 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_255_224_lpi_2,
          and_696_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_287_256 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_287_256 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_287_256_lpi_2,
          and_702_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_319_288 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_319_288 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_319_288_lpi_2,
          and_708_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_351_320 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_351_320 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_351_320_lpi_2,
          and_714_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_383_352 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_383_352 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_383_352_lpi_2,
          and_720_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_415_384 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_415_384 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_415_384_lpi_2,
          and_726_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_447_416 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_447_416 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_447_416_lpi_2,
          and_732_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_479_448 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_479_448 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_479_448_lpi_2,
          and_738_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_511_480 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_511_480 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_511_480_lpi_2,
          and_744_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_543_512 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_543_512 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_543_512_lpi_2,
          and_750_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_575_544 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_575_544 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_575_544_lpi_2,
          and_756_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_607_576 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_607_576 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_607_576_lpi_2,
          and_762_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_639_608 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_639_608 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_639_608_lpi_2,
          and_768_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_671_640 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_671_640 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_671_640_lpi_2,
          and_774_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_703_672 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_703_672 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_703_672_lpi_2,
          and_780_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_735_704 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_735_704 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_735_704_lpi_2,
          and_786_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_767_736 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_767_736 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_767_736_lpi_2,
          and_792_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_799_768 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_799_768 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_799_768_lpi_2,
          and_798_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_831_800 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_831_800 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_831_800_lpi_2,
          and_804_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_863_832 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_863_832 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_863_832_lpi_2,
          and_810_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_895_864 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_895_864 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_895_864_lpi_2,
          and_816_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_927_896 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_927_896 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_927_896_lpi_2,
          and_822_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_959_928 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_959_928 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_959_928_lpi_2,
          and_828_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_991_960 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_991_960 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_991_960_lpi_2,
          and_834_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_1023_992 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_1023_992 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1023_992_lpi_2,
          and_840_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_1055_1024 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_1055_1024 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1055_1024_lpi_2,
          and_846_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_1087_1056 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_1087_1056 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1087_1056_lpi_2,
          and_852_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_1119_1088 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_1119_1088 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1119_1088_lpi_2,
          and_858_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_1151_1120 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_1151_1120 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1151_1120_lpi_2,
          and_864_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_1183_1152 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_1183_1152 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1183_1152_lpi_2,
          and_870_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_1215_1184 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_1215_1184 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1215_1184_lpi_2,
          and_876_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_1247_1216 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_1247_1216 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1247_1216_lpi_2,
          and_882_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_1279_1248 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_1279_1248 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1279_1248_lpi_2,
          and_888_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_1311_1280 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_1311_1280 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1311_1280_lpi_2,
          and_894_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_1343_1312 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_1343_1312 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1343_1312_lpi_2,
          and_900_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_1375_1344 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_1375_1344 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1375_1344_lpi_2,
          and_906_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_1407_1376 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_1407_1376 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1407_1376_lpi_2,
          and_912_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_1439_1408 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_1439_1408 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1439_1408_lpi_2,
          and_918_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_1471_1440 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_1471_1440 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1471_1440_lpi_2,
          and_924_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_1503_1472 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_1503_1472 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1503_1472_lpi_2,
          and_930_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_1535_1504 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_1535_1504 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1535_1504_lpi_2,
          and_936_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_1567_1536 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_1567_1536 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1567_1536_lpi_2,
          and_942_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_1599_1568 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_1599_1568 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1599_1568_lpi_2,
          and_948_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_1631_1600 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_1631_1600 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1631_1600_lpi_2,
          and_954_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_1663_1632 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_1663_1632 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1663_1632_lpi_2,
          and_960_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_1695_1664 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_1695_1664 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1695_1664_lpi_2,
          and_966_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_1727_1696 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_1727_1696 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1727_1696_lpi_2,
          and_972_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_1759_1728 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_1759_1728 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1759_1728_lpi_2,
          and_978_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_1791_1760 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_1791_1760 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1791_1760_lpi_2,
          and_984_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_1823_1792 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_1823_1792 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1823_1792_lpi_2,
          and_990_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_1855_1824 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_1855_1824 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1855_1824_lpi_2,
          and_996_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_1887_1856 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_1887_1856 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1887_1856_lpi_2,
          and_1002_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_1919_1888 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_1919_1888 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1919_1888_lpi_2,
          and_1008_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_1951_1920 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_1951_1920 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1951_1920_lpi_2,
          and_1014_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_1983_1952 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_1983_1952 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_1983_1952_lpi_2,
          and_1020_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_2015_1984 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_2015_1984 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2015_1984_lpi_2,
          and_1026_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_2047_2016 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_2047_2016 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2047_2016_lpi_2,
          and_1032_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_2079_2048 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_2079_2048 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2079_2048_lpi_2,
          and_1038_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_2111_2080 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_2111_2080 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2111_2080_lpi_2,
          and_1044_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_2143_2112 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_2143_2112 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2143_2112_lpi_2,
          and_1050_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_2175_2144 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_2175_2144 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2175_2144_lpi_2,
          and_1056_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_2207_2176 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_2207_2176 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2207_2176_lpi_2,
          and_1062_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_2239_2208 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_2239_2208 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2239_2208_lpi_2,
          and_1068_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_2271_2240 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_2271_2240 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2271_2240_lpi_2,
          and_1074_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_2303_2272 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_2303_2272 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2303_2272_lpi_2,
          and_1080_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_2335_2304 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_2335_2304 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2335_2304_lpi_2,
          and_1086_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_2367_2336 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_2367_2336 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2367_2336_lpi_2,
          and_1092_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_2399_2368 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_2399_2368 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2399_2368_lpi_2,
          and_1098_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_2431_2400 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_2431_2400 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2431_2400_lpi_2,
          and_1104_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_2463_2432 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_2463_2432 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2463_2432_lpi_2,
          and_1110_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_2495_2464 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_2495_2464 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2495_2464_lpi_2,
          and_1116_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_2527_2496 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_2527_2496 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2527_2496_lpi_2,
          and_1122_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_2559_2528 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_2559_2528 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2559_2528_lpi_2,
          and_1128_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_2591_2560 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_2591_2560 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2591_2560_lpi_2,
          and_1134_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_2623_2592 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_2623_2592 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2623_2592_lpi_2,
          and_1140_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_2655_2624 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_2655_2624 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2655_2624_lpi_2,
          and_1146_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_2687_2656 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_2687_2656 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2687_2656_lpi_2,
          and_1152_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_2719_2688 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_2719_2688 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2719_2688_lpi_2,
          and_1158_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_2751_2720 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_2751_2720 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2751_2720_lpi_2,
          and_1164_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_2783_2752 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_2783_2752 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2783_2752_lpi_2,
          and_1170_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_2815_2784 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_2815_2784 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2815_2784_lpi_2,
          and_1176_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_2847_2816 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_2847_2816 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2847_2816_lpi_2,
          and_1182_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_2879_2848 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_2879_2848 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2879_2848_lpi_2,
          and_1188_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_2911_2880 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_2911_2880 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2911_2880_lpi_2,
          and_1194_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_2943_2912 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_2943_2912 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2943_2912_lpi_2,
          and_1200_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_2975_2944 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_2975_2944 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_2975_2944_lpi_2,
          and_1206_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_3007_2976 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_3007_2976 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3007_2976_lpi_2,
          and_1212_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_3039_3008 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_3039_3008 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3039_3008_lpi_2,
          and_1218_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_3071_3040 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_3071_3040 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3071_3040_lpi_2,
          and_1224_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_3103_3072 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_3103_3072 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3103_3072_lpi_2,
          and_1230_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_3135_3104 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_3135_3104 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3135_3104_lpi_2,
          and_1236_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_3167_3136 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_3167_3136 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3167_3136_lpi_2,
          and_1242_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_3199_3168 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_3199_3168 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3199_3168_lpi_2,
          and_1248_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_3231_3200 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_3231_3200 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3231_3200_lpi_2,
          and_1254_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_3263_3232 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_3263_3232 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3263_3232_lpi_2,
          and_1260_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_3295_3264 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_3295_3264 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3295_3264_lpi_2,
          and_1266_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_3327_3296 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_3327_3296 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3327_3296_lpi_2,
          and_1272_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_3359_3328 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_3359_3328 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3359_3328_lpi_2,
          and_1278_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_3391_3360 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_3391_3360 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3391_3360_lpi_2,
          and_1284_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_3423_3392 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_3423_3392 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3423_3392_lpi_2,
          and_1290_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_3455_3424 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_3455_3424 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3455_3424_lpi_2,
          and_1296_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_3487_3456 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_3487_3456 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3487_3456_lpi_2,
          and_1302_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_3519_3488 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_3519_3488 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3519_3488_lpi_2,
          and_1308_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_3551_3520 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_3551_3520 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3551_3520_lpi_2,
          and_1314_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_3583_3552 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_3583_3552 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3583_3552_lpi_2,
          and_1320_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_3615_3584 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_3615_3584 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3615_3584_lpi_2,
          and_1326_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_3647_3616 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_3647_3616 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3647_3616_lpi_2,
          and_1332_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_3679_3648 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_3679_3648 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3679_3648_lpi_2,
          and_1338_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_3711_3680 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_3711_3680 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3711_3680_lpi_2,
          and_1344_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_3743_3712 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_3743_3712 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3743_3712_lpi_2,
          and_1350_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_3775_3744 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_3775_3744 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3775_3744_lpi_2,
          and_1356_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_3807_3776 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_3807_3776 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3807_3776_lpi_2,
          and_1362_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_3839_3808 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_3839_3808 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3839_3808_lpi_2,
          and_1368_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_3871_3840 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_3871_3840 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3871_3840_lpi_2,
          and_1374_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_3903_3872 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_3903_3872 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3903_3872_lpi_2,
          and_1380_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_3935_3904 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_3935_3904 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3935_3904_lpi_2,
          and_1386_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_3967_3936 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_3967_3936 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3967_3936_lpi_2,
          and_1392_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_3999_3968 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_3999_3968 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_3999_3968_lpi_2,
          and_1398_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_4031_4000 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_4031_4000 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_4031_4000_lpi_2,
          and_1404_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_4063_4032 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_4063_4032 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_4063_4032_lpi_2,
          and_1410_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat_4095_4064 <= 32'b00000000000000000000000000000000;
    end
    else if ( fsm_output[2] ) begin
      output_rsci_idat_4095_4064 <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1, output_rsc_1_4095_4064_lpi_2,
          and_1416_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_output_rsc_triosy_obj_ld_cse <= 1'b0;
      for_equal_tmp_3 <= 1'b0;
      for_equal_tmp_5 <= 1'b0;
      for_equal_tmp_6 <= 1'b0;
      for_equal_tmp_7 <= 1'b0;
      for_equal_tmp_9 <= 1'b0;
      for_equal_tmp_10 <= 1'b0;
      for_equal_tmp_11 <= 1'b0;
      for_equal_tmp_12 <= 1'b0;
      for_equal_tmp_13 <= 1'b0;
      for_equal_tmp_14 <= 1'b0;
      for_equal_tmp_15 <= 1'b0;
      for_equal_tmp_17 <= 1'b0;
      for_equal_tmp_18 <= 1'b0;
      for_equal_tmp_19 <= 1'b0;
      for_equal_tmp_20 <= 1'b0;
      for_equal_tmp_21 <= 1'b0;
      for_equal_tmp_22 <= 1'b0;
      for_equal_tmp_23 <= 1'b0;
      for_equal_tmp_24 <= 1'b0;
      for_equal_tmp_25 <= 1'b0;
      for_equal_tmp_26 <= 1'b0;
      for_equal_tmp_27 <= 1'b0;
      for_equal_tmp_28 <= 1'b0;
      for_equal_tmp_29 <= 1'b0;
      for_equal_tmp_30 <= 1'b0;
      for_equal_tmp_31 <= 1'b0;
      for_equal_tmp_33 <= 1'b0;
      for_equal_tmp_34 <= 1'b0;
      for_equal_tmp_35 <= 1'b0;
      for_equal_tmp_36 <= 1'b0;
      for_equal_tmp_37 <= 1'b0;
      for_equal_tmp_38 <= 1'b0;
      for_equal_tmp_39 <= 1'b0;
      for_equal_tmp_40 <= 1'b0;
      for_equal_tmp_41 <= 1'b0;
      for_equal_tmp_42 <= 1'b0;
      for_equal_tmp_43 <= 1'b0;
      for_equal_tmp_44 <= 1'b0;
      for_equal_tmp_45 <= 1'b0;
      for_equal_tmp_46 <= 1'b0;
      for_equal_tmp_47 <= 1'b0;
      for_equal_tmp_48 <= 1'b0;
      for_equal_tmp_49 <= 1'b0;
      for_equal_tmp_50 <= 1'b0;
      for_equal_tmp_51 <= 1'b0;
      for_equal_tmp_52 <= 1'b0;
      for_equal_tmp_53 <= 1'b0;
      for_equal_tmp_54 <= 1'b0;
      for_equal_tmp_55 <= 1'b0;
      for_equal_tmp_56 <= 1'b0;
      for_equal_tmp_57 <= 1'b0;
      for_equal_tmp_58 <= 1'b0;
      for_equal_tmp_59 <= 1'b0;
      for_equal_tmp_60 <= 1'b0;
      for_equal_tmp_61 <= 1'b0;
      for_equal_tmp_62 <= 1'b0;
      for_equal_tmp_63 <= 1'b0;
      for_equal_tmp_65 <= 1'b0;
      for_equal_tmp_66 <= 1'b0;
      for_equal_tmp_67 <= 1'b0;
      for_equal_tmp_68 <= 1'b0;
      for_equal_tmp_69 <= 1'b0;
      for_equal_tmp_70 <= 1'b0;
      for_equal_tmp_71 <= 1'b0;
      for_equal_tmp_72 <= 1'b0;
      for_equal_tmp_73 <= 1'b0;
      for_equal_tmp_74 <= 1'b0;
      for_equal_tmp_75 <= 1'b0;
      for_equal_tmp_76 <= 1'b0;
      for_equal_tmp_77 <= 1'b0;
      for_equal_tmp_78 <= 1'b0;
      for_equal_tmp_79 <= 1'b0;
      for_equal_tmp_80 <= 1'b0;
      for_equal_tmp_81 <= 1'b0;
      for_equal_tmp_82 <= 1'b0;
      for_equal_tmp_83 <= 1'b0;
      for_equal_tmp_84 <= 1'b0;
      for_equal_tmp_85 <= 1'b0;
      for_equal_tmp_86 <= 1'b0;
      for_equal_tmp_87 <= 1'b0;
      for_equal_tmp_88 <= 1'b0;
      for_equal_tmp_89 <= 1'b0;
      for_equal_tmp_90 <= 1'b0;
      for_equal_tmp_91 <= 1'b0;
      for_equal_tmp_92 <= 1'b0;
      for_equal_tmp_93 <= 1'b0;
      for_equal_tmp_94 <= 1'b0;
      for_equal_tmp_95 <= 1'b0;
      for_equal_tmp_96 <= 1'b0;
      for_equal_tmp_97 <= 1'b0;
      for_equal_tmp_98 <= 1'b0;
      for_equal_tmp_99 <= 1'b0;
      for_equal_tmp_100 <= 1'b0;
      for_equal_tmp_101 <= 1'b0;
      for_equal_tmp_102 <= 1'b0;
      for_equal_tmp_103 <= 1'b0;
      for_equal_tmp_104 <= 1'b0;
      for_equal_tmp_105 <= 1'b0;
      for_equal_tmp_106 <= 1'b0;
      for_equal_tmp_107 <= 1'b0;
      for_equal_tmp_108 <= 1'b0;
      for_equal_tmp_109 <= 1'b0;
      for_equal_tmp_110 <= 1'b0;
      for_equal_tmp_111 <= 1'b0;
      for_equal_tmp_112 <= 1'b0;
      for_equal_tmp_113 <= 1'b0;
      for_equal_tmp_114 <= 1'b0;
      for_equal_tmp_115 <= 1'b0;
      for_equal_tmp_116 <= 1'b0;
      for_equal_tmp_117 <= 1'b0;
      for_equal_tmp_118 <= 1'b0;
      for_equal_tmp_119 <= 1'b0;
      for_equal_tmp_120 <= 1'b0;
      for_equal_tmp_121 <= 1'b0;
      for_equal_tmp_122 <= 1'b0;
      for_equal_tmp_123 <= 1'b0;
      for_equal_tmp_124 <= 1'b0;
      for_equal_tmp_125 <= 1'b0;
      for_equal_tmp_126 <= 1'b0;
      for_equal_tmp_127 <= 1'b0;
      for_nor_62_itm <= 1'b0;
      for_nor_31_itm <= 1'b0;
      for_nor_15_itm <= 1'b0;
      for_nor_7_itm <= 1'b0;
      for_nor_3_itm <= 1'b0;
      for_nor_1_itm <= 1'b0;
      for_nor_itm <= 1'b0;
      for_mux_itm <= 32'b00000000000000000000000000000000;
    end
    else begin
      reg_output_rsc_triosy_obj_ld_cse <= (i_7_0_sva_1[7]) & (fsm_output[3]);
      for_equal_tmp_3 <= (i_7_0_sva_6_0==7'b0000011);
      for_equal_tmp_5 <= (i_7_0_sva_6_0==7'b0000101);
      for_equal_tmp_6 <= (i_7_0_sva_6_0==7'b0000110);
      for_equal_tmp_7 <= (i_7_0_sva_6_0==7'b0000111);
      for_equal_tmp_9 <= (i_7_0_sva_6_0==7'b0001001);
      for_equal_tmp_10 <= (i_7_0_sva_6_0==7'b0001010);
      for_equal_tmp_11 <= (i_7_0_sva_6_0==7'b0001011);
      for_equal_tmp_12 <= (i_7_0_sva_6_0==7'b0001100);
      for_equal_tmp_13 <= (i_7_0_sva_6_0==7'b0001101);
      for_equal_tmp_14 <= (i_7_0_sva_6_0==7'b0001110);
      for_equal_tmp_15 <= (i_7_0_sva_6_0==7'b0001111);
      for_equal_tmp_17 <= (i_7_0_sva_6_0==7'b0010001);
      for_equal_tmp_18 <= (i_7_0_sva_6_0==7'b0010010);
      for_equal_tmp_19 <= (i_7_0_sva_6_0==7'b0010011);
      for_equal_tmp_20 <= (i_7_0_sva_6_0==7'b0010100);
      for_equal_tmp_21 <= (i_7_0_sva_6_0==7'b0010101);
      for_equal_tmp_22 <= (i_7_0_sva_6_0==7'b0010110);
      for_equal_tmp_23 <= (i_7_0_sva_6_0==7'b0010111);
      for_equal_tmp_24 <= (i_7_0_sva_6_0==7'b0011000);
      for_equal_tmp_25 <= (i_7_0_sva_6_0==7'b0011001);
      for_equal_tmp_26 <= (i_7_0_sva_6_0==7'b0011010);
      for_equal_tmp_27 <= (i_7_0_sva_6_0==7'b0011011);
      for_equal_tmp_28 <= (i_7_0_sva_6_0==7'b0011100);
      for_equal_tmp_29 <= (i_7_0_sva_6_0==7'b0011101);
      for_equal_tmp_30 <= (i_7_0_sva_6_0==7'b0011110);
      for_equal_tmp_31 <= (i_7_0_sva_6_0==7'b0011111);
      for_equal_tmp_33 <= (i_7_0_sva_6_0==7'b0100001);
      for_equal_tmp_34 <= (i_7_0_sva_6_0==7'b0100010);
      for_equal_tmp_35 <= (i_7_0_sva_6_0==7'b0100011);
      for_equal_tmp_36 <= (i_7_0_sva_6_0==7'b0100100);
      for_equal_tmp_37 <= (i_7_0_sva_6_0==7'b0100101);
      for_equal_tmp_38 <= (i_7_0_sva_6_0==7'b0100110);
      for_equal_tmp_39 <= (i_7_0_sva_6_0==7'b0100111);
      for_equal_tmp_40 <= (i_7_0_sva_6_0==7'b0101000);
      for_equal_tmp_41 <= (i_7_0_sva_6_0==7'b0101001);
      for_equal_tmp_42 <= (i_7_0_sva_6_0==7'b0101010);
      for_equal_tmp_43 <= (i_7_0_sva_6_0==7'b0101011);
      for_equal_tmp_44 <= (i_7_0_sva_6_0==7'b0101100);
      for_equal_tmp_45 <= (i_7_0_sva_6_0==7'b0101101);
      for_equal_tmp_46 <= (i_7_0_sva_6_0==7'b0101110);
      for_equal_tmp_47 <= (i_7_0_sva_6_0==7'b0101111);
      for_equal_tmp_48 <= (i_7_0_sva_6_0==7'b0110000);
      for_equal_tmp_49 <= (i_7_0_sva_6_0==7'b0110001);
      for_equal_tmp_50 <= (i_7_0_sva_6_0==7'b0110010);
      for_equal_tmp_51 <= (i_7_0_sva_6_0==7'b0110011);
      for_equal_tmp_52 <= (i_7_0_sva_6_0==7'b0110100);
      for_equal_tmp_53 <= (i_7_0_sva_6_0==7'b0110101);
      for_equal_tmp_54 <= (i_7_0_sva_6_0==7'b0110110);
      for_equal_tmp_55 <= (i_7_0_sva_6_0==7'b0110111);
      for_equal_tmp_56 <= (i_7_0_sva_6_0==7'b0111000);
      for_equal_tmp_57 <= (i_7_0_sva_6_0==7'b0111001);
      for_equal_tmp_58 <= (i_7_0_sva_6_0==7'b0111010);
      for_equal_tmp_59 <= (i_7_0_sva_6_0==7'b0111011);
      for_equal_tmp_60 <= (i_7_0_sva_6_0==7'b0111100);
      for_equal_tmp_61 <= (i_7_0_sva_6_0==7'b0111101);
      for_equal_tmp_62 <= (i_7_0_sva_6_0==7'b0111110);
      for_equal_tmp_63 <= (i_7_0_sva_6_0==7'b0111111);
      for_equal_tmp_65 <= (i_7_0_sva_6_0==7'b1000001);
      for_equal_tmp_66 <= (i_7_0_sva_6_0==7'b1000010);
      for_equal_tmp_67 <= (i_7_0_sva_6_0==7'b1000011);
      for_equal_tmp_68 <= (i_7_0_sva_6_0==7'b1000100);
      for_equal_tmp_69 <= (i_7_0_sva_6_0==7'b1000101);
      for_equal_tmp_70 <= (i_7_0_sva_6_0==7'b1000110);
      for_equal_tmp_71 <= (i_7_0_sva_6_0==7'b1000111);
      for_equal_tmp_72 <= (i_7_0_sva_6_0==7'b1001000);
      for_equal_tmp_73 <= (i_7_0_sva_6_0==7'b1001001);
      for_equal_tmp_74 <= (i_7_0_sva_6_0==7'b1001010);
      for_equal_tmp_75 <= (i_7_0_sva_6_0==7'b1001011);
      for_equal_tmp_76 <= (i_7_0_sva_6_0==7'b1001100);
      for_equal_tmp_77 <= (i_7_0_sva_6_0==7'b1001101);
      for_equal_tmp_78 <= (i_7_0_sva_6_0==7'b1001110);
      for_equal_tmp_79 <= (i_7_0_sva_6_0==7'b1001111);
      for_equal_tmp_80 <= (i_7_0_sva_6_0==7'b1010000);
      for_equal_tmp_81 <= (i_7_0_sva_6_0==7'b1010001);
      for_equal_tmp_82 <= (i_7_0_sva_6_0==7'b1010010);
      for_equal_tmp_83 <= (i_7_0_sva_6_0==7'b1010011);
      for_equal_tmp_84 <= (i_7_0_sva_6_0==7'b1010100);
      for_equal_tmp_85 <= (i_7_0_sva_6_0==7'b1010101);
      for_equal_tmp_86 <= (i_7_0_sva_6_0==7'b1010110);
      for_equal_tmp_87 <= (i_7_0_sva_6_0==7'b1010111);
      for_equal_tmp_88 <= (i_7_0_sva_6_0==7'b1011000);
      for_equal_tmp_89 <= (i_7_0_sva_6_0==7'b1011001);
      for_equal_tmp_90 <= (i_7_0_sva_6_0==7'b1011010);
      for_equal_tmp_91 <= (i_7_0_sva_6_0==7'b1011011);
      for_equal_tmp_92 <= (i_7_0_sva_6_0==7'b1011100);
      for_equal_tmp_93 <= (i_7_0_sva_6_0==7'b1011101);
      for_equal_tmp_94 <= (i_7_0_sva_6_0==7'b1011110);
      for_equal_tmp_95 <= (i_7_0_sva_6_0==7'b1011111);
      for_equal_tmp_96 <= (i_7_0_sva_6_0==7'b1100000);
      for_equal_tmp_97 <= (i_7_0_sva_6_0==7'b1100001);
      for_equal_tmp_98 <= (i_7_0_sva_6_0==7'b1100010);
      for_equal_tmp_99 <= (i_7_0_sva_6_0==7'b1100011);
      for_equal_tmp_100 <= (i_7_0_sva_6_0==7'b1100100);
      for_equal_tmp_101 <= (i_7_0_sva_6_0==7'b1100101);
      for_equal_tmp_102 <= (i_7_0_sva_6_0==7'b1100110);
      for_equal_tmp_103 <= (i_7_0_sva_6_0==7'b1100111);
      for_equal_tmp_104 <= (i_7_0_sva_6_0==7'b1101000);
      for_equal_tmp_105 <= (i_7_0_sva_6_0==7'b1101001);
      for_equal_tmp_106 <= (i_7_0_sva_6_0==7'b1101010);
      for_equal_tmp_107 <= (i_7_0_sva_6_0==7'b1101011);
      for_equal_tmp_108 <= (i_7_0_sva_6_0==7'b1101100);
      for_equal_tmp_109 <= (i_7_0_sva_6_0==7'b1101101);
      for_equal_tmp_110 <= (i_7_0_sva_6_0==7'b1101110);
      for_equal_tmp_111 <= (i_7_0_sva_6_0==7'b1101111);
      for_equal_tmp_112 <= (i_7_0_sva_6_0==7'b1110000);
      for_equal_tmp_113 <= (i_7_0_sva_6_0==7'b1110001);
      for_equal_tmp_114 <= (i_7_0_sva_6_0==7'b1110010);
      for_equal_tmp_115 <= (i_7_0_sva_6_0==7'b1110011);
      for_equal_tmp_116 <= (i_7_0_sva_6_0==7'b1110100);
      for_equal_tmp_117 <= (i_7_0_sva_6_0==7'b1110101);
      for_equal_tmp_118 <= (i_7_0_sva_6_0==7'b1110110);
      for_equal_tmp_119 <= (i_7_0_sva_6_0==7'b1110111);
      for_equal_tmp_120 <= (i_7_0_sva_6_0==7'b1111000);
      for_equal_tmp_121 <= (i_7_0_sva_6_0==7'b1111001);
      for_equal_tmp_122 <= (i_7_0_sva_6_0==7'b1111010);
      for_equal_tmp_123 <= (i_7_0_sva_6_0==7'b1111011);
      for_equal_tmp_124 <= (i_7_0_sva_6_0==7'b1111100);
      for_equal_tmp_125 <= (i_7_0_sva_6_0==7'b1111101);
      for_equal_tmp_126 <= (i_7_0_sva_6_0==7'b1111110);
      for_equal_tmp_127 <= (i_7_0_sva_6_0==7'b1111111);
      for_nor_62_itm <= ~((i_7_0_sva_6_0[5:0]!=6'b000000));
      for_nor_31_itm <= ~((i_7_0_sva_6_0[6]) | (i_7_0_sva_6_0[4]) | (i_7_0_sva_6_0[3])
          | (i_7_0_sva_6_0[2]) | (i_7_0_sva_6_0[1]) | (i_7_0_sva_6_0[0]));
      for_nor_15_itm <= ~((i_7_0_sva_6_0[6]) | (i_7_0_sva_6_0[5]) | (i_7_0_sva_6_0[3])
          | (i_7_0_sva_6_0[2]) | (i_7_0_sva_6_0[1]) | (i_7_0_sva_6_0[0]));
      for_nor_7_itm <= ~((i_7_0_sva_6_0[6]) | (i_7_0_sva_6_0[5]) | (i_7_0_sva_6_0[4])
          | (i_7_0_sva_6_0[2]) | (i_7_0_sva_6_0[1]) | (i_7_0_sva_6_0[0]));
      for_nor_3_itm <= ~((i_7_0_sva_6_0[6]) | (i_7_0_sva_6_0[5]) | (i_7_0_sva_6_0[4])
          | (i_7_0_sva_6_0[3]) | (i_7_0_sva_6_0[1]) | (i_7_0_sva_6_0[0]));
      for_nor_1_itm <= ~((i_7_0_sva_6_0[6]) | (i_7_0_sva_6_0[5]) | (i_7_0_sva_6_0[4])
          | (i_7_0_sva_6_0[3]) | (i_7_0_sva_6_0[2]) | (i_7_0_sva_6_0[0]));
      for_nor_itm <= ~((i_7_0_sva_6_0[6:1]!=6'b000000));
      for_mux_itm <= MUX_v_32_128_2((input_rsci_idat[31:0]), (input_rsci_idat[63:32]),
          (input_rsci_idat[95:64]), (input_rsci_idat[127:96]), (input_rsci_idat[159:128]),
          (input_rsci_idat[191:160]), (input_rsci_idat[223:192]), (input_rsci_idat[255:224]),
          (input_rsci_idat[287:256]), (input_rsci_idat[319:288]), (input_rsci_idat[351:320]),
          (input_rsci_idat[383:352]), (input_rsci_idat[415:384]), (input_rsci_idat[447:416]),
          (input_rsci_idat[479:448]), (input_rsci_idat[511:480]), (input_rsci_idat[543:512]),
          (input_rsci_idat[575:544]), (input_rsci_idat[607:576]), (input_rsci_idat[639:608]),
          (input_rsci_idat[671:640]), (input_rsci_idat[703:672]), (input_rsci_idat[735:704]),
          (input_rsci_idat[767:736]), (input_rsci_idat[799:768]), (input_rsci_idat[831:800]),
          (input_rsci_idat[863:832]), (input_rsci_idat[895:864]), (input_rsci_idat[927:896]),
          (input_rsci_idat[959:928]), (input_rsci_idat[991:960]), (input_rsci_idat[1023:992]),
          (input_rsci_idat[1055:1024]), (input_rsci_idat[1087:1056]), (input_rsci_idat[1119:1088]),
          (input_rsci_idat[1151:1120]), (input_rsci_idat[1183:1152]), (input_rsci_idat[1215:1184]),
          (input_rsci_idat[1247:1216]), (input_rsci_idat[1279:1248]), (input_rsci_idat[1311:1280]),
          (input_rsci_idat[1343:1312]), (input_rsci_idat[1375:1344]), (input_rsci_idat[1407:1376]),
          (input_rsci_idat[1439:1408]), (input_rsci_idat[1471:1440]), (input_rsci_idat[1503:1472]),
          (input_rsci_idat[1535:1504]), (input_rsci_idat[1567:1536]), (input_rsci_idat[1599:1568]),
          (input_rsci_idat[1631:1600]), (input_rsci_idat[1663:1632]), (input_rsci_idat[1695:1664]),
          (input_rsci_idat[1727:1696]), (input_rsci_idat[1759:1728]), (input_rsci_idat[1791:1760]),
          (input_rsci_idat[1823:1792]), (input_rsci_idat[1855:1824]), (input_rsci_idat[1887:1856]),
          (input_rsci_idat[1919:1888]), (input_rsci_idat[1951:1920]), (input_rsci_idat[1983:1952]),
          (input_rsci_idat[2015:1984]), (input_rsci_idat[2047:2016]), (input_rsci_idat[2079:2048]),
          (input_rsci_idat[2111:2080]), (input_rsci_idat[2143:2112]), (input_rsci_idat[2175:2144]),
          (input_rsci_idat[2207:2176]), (input_rsci_idat[2239:2208]), (input_rsci_idat[2271:2240]),
          (input_rsci_idat[2303:2272]), (input_rsci_idat[2335:2304]), (input_rsci_idat[2367:2336]),
          (input_rsci_idat[2399:2368]), (input_rsci_idat[2431:2400]), (input_rsci_idat[2463:2432]),
          (input_rsci_idat[2495:2464]), (input_rsci_idat[2527:2496]), (input_rsci_idat[2559:2528]),
          (input_rsci_idat[2591:2560]), (input_rsci_idat[2623:2592]), (input_rsci_idat[2655:2624]),
          (input_rsci_idat[2687:2656]), (input_rsci_idat[2719:2688]), (input_rsci_idat[2751:2720]),
          (input_rsci_idat[2783:2752]), (input_rsci_idat[2815:2784]), (input_rsci_idat[2847:2816]),
          (input_rsci_idat[2879:2848]), (input_rsci_idat[2911:2880]), (input_rsci_idat[2943:2912]),
          (input_rsci_idat[2975:2944]), (input_rsci_idat[3007:2976]), (input_rsci_idat[3039:3008]),
          (input_rsci_idat[3071:3040]), (input_rsci_idat[3103:3072]), (input_rsci_idat[3135:3104]),
          (input_rsci_idat[3167:3136]), (input_rsci_idat[3199:3168]), (input_rsci_idat[3231:3200]),
          (input_rsci_idat[3263:3232]), (input_rsci_idat[3295:3264]), (input_rsci_idat[3327:3296]),
          (input_rsci_idat[3359:3328]), (input_rsci_idat[3391:3360]), (input_rsci_idat[3423:3392]),
          (input_rsci_idat[3455:3424]), (input_rsci_idat[3487:3456]), (input_rsci_idat[3519:3488]),
          (input_rsci_idat[3551:3520]), (input_rsci_idat[3583:3552]), (input_rsci_idat[3615:3584]),
          (input_rsci_idat[3647:3616]), (input_rsci_idat[3679:3648]), (input_rsci_idat[3711:3680]),
          (input_rsci_idat[3743:3712]), (input_rsci_idat[3775:3744]), (input_rsci_idat[3807:3776]),
          (input_rsci_idat[3839:3808]), (input_rsci_idat[3871:3840]), (input_rsci_idat[3903:3872]),
          (input_rsci_idat[3935:3904]), (input_rsci_idat[3967:3936]), (input_rsci_idat[3999:3968]),
          (input_rsci_idat[4031:4000]), (input_rsci_idat[4063:4032]), (input_rsci_idat[4095:4064]),
          i_7_0_sva_6_0);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_2047_2016_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_2047_2016_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2047_2016_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_253_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_2079_2048_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_2079_2048_lpi_2_dfm <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1,
          output_rsc_1_2079_2048_lpi_2, for_and_251_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_2015_1984_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_2015_1984_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2015_1984_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_249_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_2111_2080_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_2111_2080_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2111_2080_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_247_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_1983_1952_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_1983_1952_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1983_1952_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_245_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_2143_2112_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_2143_2112_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2143_2112_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_243_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_1951_1920_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_1951_1920_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1951_1920_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_241_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_2175_2144_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_2175_2144_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2175_2144_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_239_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_1919_1888_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_1919_1888_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1919_1888_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_237_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_2207_2176_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_2207_2176_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2207_2176_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_235_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_1887_1856_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_1887_1856_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1887_1856_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_233_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_2239_2208_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_2239_2208_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2239_2208_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_231_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_1855_1824_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_1855_1824_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1855_1824_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_229_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_2271_2240_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_2271_2240_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2271_2240_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_227_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_1823_1792_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_1823_1792_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1823_1792_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_225_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_2303_2272_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_2303_2272_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2303_2272_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_223_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_1791_1760_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_1791_1760_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1791_1760_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_221_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_2335_2304_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_2335_2304_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2335_2304_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_219_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_1759_1728_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_1759_1728_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1759_1728_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_217_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_2367_2336_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_2367_2336_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2367_2336_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_215_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_1727_1696_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_1727_1696_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1727_1696_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_213_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_2399_2368_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_2399_2368_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2399_2368_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_211_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_1695_1664_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_1695_1664_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1695_1664_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_209_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_2431_2400_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_2431_2400_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2431_2400_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_207_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_1663_1632_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_1663_1632_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1663_1632_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_205_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_2463_2432_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_2463_2432_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2463_2432_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_203_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_1631_1600_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_1631_1600_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1631_1600_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_201_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_2495_2464_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_2495_2464_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2495_2464_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_199_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_1599_1568_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_1599_1568_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1599_1568_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_197_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_2527_2496_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_2527_2496_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2527_2496_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_195_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_1567_1536_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_1567_1536_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1567_1536_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_193_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_2559_2528_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_2559_2528_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2559_2528_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_191_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_1535_1504_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_1535_1504_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1535_1504_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_189_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_2591_2560_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_2591_2560_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2591_2560_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_187_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_1503_1472_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_1503_1472_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1503_1472_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_185_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_2623_2592_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_2623_2592_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2623_2592_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_183_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_1471_1440_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_1471_1440_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1471_1440_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_181_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_2655_2624_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_2655_2624_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2655_2624_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_179_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_1439_1408_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_1439_1408_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1439_1408_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_177_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_2687_2656_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_2687_2656_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2687_2656_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_175_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_1407_1376_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_1407_1376_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1407_1376_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_173_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_2719_2688_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_2719_2688_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2719_2688_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_171_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_1375_1344_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_1375_1344_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1375_1344_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_169_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_2751_2720_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_2751_2720_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2751_2720_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_167_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_1343_1312_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_1343_1312_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1343_1312_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_165_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_2783_2752_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_2783_2752_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2783_2752_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_163_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_1311_1280_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_1311_1280_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1311_1280_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_161_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_2815_2784_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_2815_2784_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2815_2784_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_159_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_1279_1248_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_1279_1248_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1279_1248_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_157_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_2847_2816_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_2847_2816_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2847_2816_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_155_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_1247_1216_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_1247_1216_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1247_1216_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_153_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_2879_2848_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_2879_2848_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2879_2848_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_151_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_1215_1184_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_1215_1184_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1215_1184_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_149_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_2911_2880_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_2911_2880_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2911_2880_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_147_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_1183_1152_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_1183_1152_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1183_1152_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_145_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_2943_2912_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_2943_2912_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2943_2912_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_143_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_1151_1120_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_1151_1120_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1151_1120_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_141_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_2975_2944_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_2975_2944_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_2975_2944_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_139_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_1119_1088_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_1119_1088_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1119_1088_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_137_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_3007_2976_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_3007_2976_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3007_2976_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_135_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_1087_1056_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_1087_1056_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1087_1056_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_133_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_3039_3008_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_3039_3008_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3039_3008_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_131_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_1055_1024_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_1055_1024_lpi_2_dfm <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1,
          output_rsc_1_1055_1024_lpi_2, for_and_129_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_3071_3040_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_3071_3040_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3071_3040_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_127_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_1023_992_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_1023_992_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_1023_992_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_125_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_3103_3072_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_3103_3072_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3103_3072_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_123_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_991_960_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_991_960_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_991_960_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_121_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_3135_3104_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_3135_3104_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3135_3104_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_119_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_959_928_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_959_928_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_959_928_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_117_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_3167_3136_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_3167_3136_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3167_3136_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_115_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_927_896_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_927_896_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_927_896_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_113_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_3199_3168_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_3199_3168_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3199_3168_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_111_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_895_864_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_895_864_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_895_864_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_109_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_3231_3200_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_3231_3200_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3231_3200_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_107_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_863_832_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_863_832_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_863_832_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_105_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_3263_3232_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_3263_3232_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3263_3232_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_103_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_831_800_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_831_800_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_831_800_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_101_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_3295_3264_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_3295_3264_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3295_3264_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_99_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_799_768_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_799_768_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_799_768_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_97_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_3327_3296_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_3327_3296_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3327_3296_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_95_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_767_736_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_767_736_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_767_736_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_93_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_3359_3328_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_3359_3328_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3359_3328_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_91_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_735_704_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_735_704_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_735_704_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_89_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_3391_3360_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_3391_3360_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3391_3360_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_87_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_703_672_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_703_672_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_703_672_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_85_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_3423_3392_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_3423_3392_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3423_3392_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_83_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_671_640_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_671_640_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_671_640_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_81_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_3455_3424_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_3455_3424_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3455_3424_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_79_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_639_608_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_639_608_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_639_608_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_77_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_3487_3456_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_3487_3456_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3487_3456_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_75_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_607_576_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_607_576_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_607_576_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_73_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_3519_3488_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_3519_3488_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3519_3488_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_71_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_575_544_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_575_544_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_575_544_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_69_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_3551_3520_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_3551_3520_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3551_3520_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_67_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_543_512_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_543_512_lpi_2_dfm <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1,
          output_rsc_1_543_512_lpi_2, for_and_65_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_3583_3552_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_3583_3552_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3583_3552_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_63_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_511_480_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_511_480_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_511_480_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_61_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_3615_3584_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_3615_3584_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3615_3584_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_59_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_479_448_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_479_448_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_479_448_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_57_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_3647_3616_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_3647_3616_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3647_3616_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_55_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_447_416_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_447_416_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_447_416_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_53_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_3679_3648_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_3679_3648_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3679_3648_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_51_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_415_384_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_415_384_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_415_384_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_49_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_3711_3680_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_3711_3680_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3711_3680_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_47_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_383_352_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_383_352_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_383_352_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_45_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_3743_3712_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_3743_3712_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3743_3712_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_43_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_351_320_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_351_320_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_351_320_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_41_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_3775_3744_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_3775_3744_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3775_3744_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_39_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_319_288_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_319_288_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_319_288_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_37_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_3807_3776_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_3807_3776_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3807_3776_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_35_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_287_256_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_287_256_lpi_2_dfm <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1,
          output_rsc_1_287_256_lpi_2, for_and_33_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_3839_3808_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_3839_3808_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3839_3808_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_31_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_255_224_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_255_224_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_255_224_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_29_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_3871_3840_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_3871_3840_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3871_3840_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_27_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_223_192_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_223_192_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_223_192_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_25_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_3903_3872_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_3903_3872_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3903_3872_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_23_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_191_160_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_191_160_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_191_160_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_21_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_3935_3904_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_3935_3904_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3935_3904_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_19_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_159_128_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_159_128_lpi_2_dfm <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1,
          output_rsc_1_159_128_lpi_2, for_and_17_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_3967_3936_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_3967_3936_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3967_3936_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_15_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_127_96_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_127_96_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_127_96_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_13_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_3999_3968_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_3999_3968_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_3999_3968_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_11_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_95_64_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_95_64_lpi_2_dfm <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1,
          output_rsc_1_95_64_lpi_2, for_and_9_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_4031_4000_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_4031_4000_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_4031_4000_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_7_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_63_32_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_63_32_lpi_2_dfm <= MUX_v_32_2_2(for_for_mul_1_cmx_sva_1,
          output_rsc_1_63_32_lpi_2, for_and_5_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_4063_4032_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_4063_4032_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_4063_4032_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_3_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_31_0_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_31_0_lpi_2_dfm <= output_output_mux_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_io_read_output_rsc_sdt_4095_4064_lpi_2_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_tmp_643 ) begin
      for_io_read_output_rsc_sdt_4095_4064_lpi_2_dfm <= MUX_v_32_2_2(output_rsc_1_4095_4064_lpi_2,
          for_for_mul_1_cmx_sva_1, for_and_1_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      i_7_0_sva_1 <= 8'b00000000;
    end
    else if ( fsm_output[1] ) begin
      i_7_0_sva_1 <= nl_i_7_0_sva_1[7:0];
    end
  end
  assign and_660_nl = or_dcpl_330 & (fsm_output[2]);
  assign and_666_nl = or_dcpl_331 & (fsm_output[2]);
  assign and_672_nl = (~ for_equal_tmp_3) & (fsm_output[2]);
  assign and_678_nl = or_dcpl_332 & (fsm_output[2]);
  assign and_684_nl = (~ for_equal_tmp_5) & (fsm_output[2]);
  assign and_690_nl = (~ for_equal_tmp_6) & (fsm_output[2]);
  assign and_696_nl = (~ for_equal_tmp_7) & (fsm_output[2]);
  assign and_702_nl = or_dcpl_333 & (fsm_output[2]);
  assign and_708_nl = (~ for_equal_tmp_9) & (fsm_output[2]);
  assign and_714_nl = (~ for_equal_tmp_10) & (fsm_output[2]);
  assign and_720_nl = (~ for_equal_tmp_11) & (fsm_output[2]);
  assign and_726_nl = (~ for_equal_tmp_12) & (fsm_output[2]);
  assign and_732_nl = (~ for_equal_tmp_13) & (fsm_output[2]);
  assign and_738_nl = (~ for_equal_tmp_14) & (fsm_output[2]);
  assign and_744_nl = (~ for_equal_tmp_15) & (fsm_output[2]);
  assign and_750_nl = or_dcpl_334 & (fsm_output[2]);
  assign and_756_nl = (~ for_equal_tmp_17) & (fsm_output[2]);
  assign and_762_nl = (~ for_equal_tmp_18) & (fsm_output[2]);
  assign and_768_nl = (~ for_equal_tmp_19) & (fsm_output[2]);
  assign and_774_nl = (~ for_equal_tmp_20) & (fsm_output[2]);
  assign and_780_nl = (~ for_equal_tmp_21) & (fsm_output[2]);
  assign and_786_nl = (~ for_equal_tmp_22) & (fsm_output[2]);
  assign and_792_nl = (~ for_equal_tmp_23) & (fsm_output[2]);
  assign and_798_nl = (~ for_equal_tmp_24) & (fsm_output[2]);
  assign and_804_nl = (~ for_equal_tmp_25) & (fsm_output[2]);
  assign and_810_nl = (~ for_equal_tmp_26) & (fsm_output[2]);
  assign and_816_nl = (~ for_equal_tmp_27) & (fsm_output[2]);
  assign and_822_nl = (~ for_equal_tmp_28) & (fsm_output[2]);
  assign and_828_nl = (~ for_equal_tmp_29) & (fsm_output[2]);
  assign and_834_nl = (~ for_equal_tmp_30) & (fsm_output[2]);
  assign and_840_nl = (~ for_equal_tmp_31) & (fsm_output[2]);
  assign and_846_nl = or_dcpl_335 & (fsm_output[2]);
  assign and_852_nl = (~ for_equal_tmp_33) & (fsm_output[2]);
  assign and_858_nl = (~ for_equal_tmp_34) & (fsm_output[2]);
  assign and_864_nl = (~ for_equal_tmp_35) & (fsm_output[2]);
  assign and_870_nl = (~ for_equal_tmp_36) & (fsm_output[2]);
  assign and_876_nl = (~ for_equal_tmp_37) & (fsm_output[2]);
  assign and_882_nl = (~ for_equal_tmp_38) & (fsm_output[2]);
  assign and_888_nl = (~ for_equal_tmp_39) & (fsm_output[2]);
  assign and_894_nl = (~ for_equal_tmp_40) & (fsm_output[2]);
  assign and_900_nl = (~ for_equal_tmp_41) & (fsm_output[2]);
  assign and_906_nl = (~ for_equal_tmp_42) & (fsm_output[2]);
  assign and_912_nl = (~ for_equal_tmp_43) & (fsm_output[2]);
  assign and_918_nl = (~ for_equal_tmp_44) & (fsm_output[2]);
  assign and_924_nl = (~ for_equal_tmp_45) & (fsm_output[2]);
  assign and_930_nl = (~ for_equal_tmp_46) & (fsm_output[2]);
  assign and_936_nl = (~ for_equal_tmp_47) & (fsm_output[2]);
  assign and_942_nl = (~ for_equal_tmp_48) & (fsm_output[2]);
  assign and_948_nl = (~ for_equal_tmp_49) & (fsm_output[2]);
  assign and_954_nl = (~ for_equal_tmp_50) & (fsm_output[2]);
  assign and_960_nl = (~ for_equal_tmp_51) & (fsm_output[2]);
  assign and_966_nl = (~ for_equal_tmp_52) & (fsm_output[2]);
  assign and_972_nl = (~ for_equal_tmp_53) & (fsm_output[2]);
  assign and_978_nl = (~ for_equal_tmp_54) & (fsm_output[2]);
  assign and_984_nl = (~ for_equal_tmp_55) & (fsm_output[2]);
  assign and_990_nl = (~ for_equal_tmp_56) & (fsm_output[2]);
  assign and_996_nl = (~ for_equal_tmp_57) & (fsm_output[2]);
  assign and_1002_nl = (~ for_equal_tmp_58) & (fsm_output[2]);
  assign and_1008_nl = (~ for_equal_tmp_59) & (fsm_output[2]);
  assign and_1014_nl = (~ for_equal_tmp_60) & (fsm_output[2]);
  assign and_1020_nl = (~ for_equal_tmp_61) & (fsm_output[2]);
  assign and_1026_nl = (~ for_equal_tmp_62) & (fsm_output[2]);
  assign and_1032_nl = (~ for_equal_tmp_63) & (fsm_output[2]);
  assign and_1038_nl = or_dcpl_336 & (fsm_output[2]);
  assign and_1044_nl = (~ for_equal_tmp_65) & (fsm_output[2]);
  assign and_1050_nl = (~ for_equal_tmp_66) & (fsm_output[2]);
  assign and_1056_nl = (~ for_equal_tmp_67) & (fsm_output[2]);
  assign and_1062_nl = (~ for_equal_tmp_68) & (fsm_output[2]);
  assign and_1068_nl = (~ for_equal_tmp_69) & (fsm_output[2]);
  assign and_1074_nl = (~ for_equal_tmp_70) & (fsm_output[2]);
  assign and_1080_nl = (~ for_equal_tmp_71) & (fsm_output[2]);
  assign and_1086_nl = (~ for_equal_tmp_72) & (fsm_output[2]);
  assign and_1092_nl = (~ for_equal_tmp_73) & (fsm_output[2]);
  assign and_1098_nl = (~ for_equal_tmp_74) & (fsm_output[2]);
  assign and_1104_nl = (~ for_equal_tmp_75) & (fsm_output[2]);
  assign and_1110_nl = (~ for_equal_tmp_76) & (fsm_output[2]);
  assign and_1116_nl = (~ for_equal_tmp_77) & (fsm_output[2]);
  assign and_1122_nl = (~ for_equal_tmp_78) & (fsm_output[2]);
  assign and_1128_nl = (~ for_equal_tmp_79) & (fsm_output[2]);
  assign and_1134_nl = (~ for_equal_tmp_80) & (fsm_output[2]);
  assign and_1140_nl = (~ for_equal_tmp_81) & (fsm_output[2]);
  assign and_1146_nl = (~ for_equal_tmp_82) & (fsm_output[2]);
  assign and_1152_nl = (~ for_equal_tmp_83) & (fsm_output[2]);
  assign and_1158_nl = (~ for_equal_tmp_84) & (fsm_output[2]);
  assign and_1164_nl = (~ for_equal_tmp_85) & (fsm_output[2]);
  assign and_1170_nl = (~ for_equal_tmp_86) & (fsm_output[2]);
  assign and_1176_nl = (~ for_equal_tmp_87) & (fsm_output[2]);
  assign and_1182_nl = (~ for_equal_tmp_88) & (fsm_output[2]);
  assign and_1188_nl = (~ for_equal_tmp_89) & (fsm_output[2]);
  assign and_1194_nl = (~ for_equal_tmp_90) & (fsm_output[2]);
  assign and_1200_nl = (~ for_equal_tmp_91) & (fsm_output[2]);
  assign and_1206_nl = (~ for_equal_tmp_92) & (fsm_output[2]);
  assign and_1212_nl = (~ for_equal_tmp_93) & (fsm_output[2]);
  assign and_1218_nl = (~ for_equal_tmp_94) & (fsm_output[2]);
  assign and_1224_nl = (~ for_equal_tmp_95) & (fsm_output[2]);
  assign and_1230_nl = (~ for_equal_tmp_96) & (fsm_output[2]);
  assign and_1236_nl = (~ for_equal_tmp_97) & (fsm_output[2]);
  assign and_1242_nl = (~ for_equal_tmp_98) & (fsm_output[2]);
  assign and_1248_nl = (~ for_equal_tmp_99) & (fsm_output[2]);
  assign and_1254_nl = (~ for_equal_tmp_100) & (fsm_output[2]);
  assign and_1260_nl = (~ for_equal_tmp_101) & (fsm_output[2]);
  assign and_1266_nl = (~ for_equal_tmp_102) & (fsm_output[2]);
  assign and_1272_nl = (~ for_equal_tmp_103) & (fsm_output[2]);
  assign and_1278_nl = (~ for_equal_tmp_104) & (fsm_output[2]);
  assign and_1284_nl = (~ for_equal_tmp_105) & (fsm_output[2]);
  assign and_1290_nl = (~ for_equal_tmp_106) & (fsm_output[2]);
  assign and_1296_nl = (~ for_equal_tmp_107) & (fsm_output[2]);
  assign and_1302_nl = (~ for_equal_tmp_108) & (fsm_output[2]);
  assign and_1308_nl = (~ for_equal_tmp_109) & (fsm_output[2]);
  assign and_1314_nl = (~ for_equal_tmp_110) & (fsm_output[2]);
  assign and_1320_nl = (~ for_equal_tmp_111) & (fsm_output[2]);
  assign and_1326_nl = (~ for_equal_tmp_112) & (fsm_output[2]);
  assign and_1332_nl = (~ for_equal_tmp_113) & (fsm_output[2]);
  assign and_1338_nl = (~ for_equal_tmp_114) & (fsm_output[2]);
  assign and_1344_nl = (~ for_equal_tmp_115) & (fsm_output[2]);
  assign and_1350_nl = (~ for_equal_tmp_116) & (fsm_output[2]);
  assign and_1356_nl = (~ for_equal_tmp_117) & (fsm_output[2]);
  assign and_1362_nl = (~ for_equal_tmp_118) & (fsm_output[2]);
  assign and_1368_nl = (~ for_equal_tmp_119) & (fsm_output[2]);
  assign and_1374_nl = (~ for_equal_tmp_120) & (fsm_output[2]);
  assign and_1380_nl = (~ for_equal_tmp_121) & (fsm_output[2]);
  assign and_1386_nl = (~ for_equal_tmp_122) & (fsm_output[2]);
  assign and_1392_nl = (~ for_equal_tmp_123) & (fsm_output[2]);
  assign and_1398_nl = (~ for_equal_tmp_124) & (fsm_output[2]);
  assign and_1404_nl = (~ for_equal_tmp_125) & (fsm_output[2]);
  assign and_1410_nl = (~ for_equal_tmp_126) & (fsm_output[2]);
  assign and_1416_nl = (~ for_equal_tmp_127) & (fsm_output[2]);
  assign for_and_253_nl = for_equal_tmp_63 & (~ or_tmp_643);
  assign for_and_251_nl = or_dcpl_336 & (~ or_tmp_643);
  assign for_and_249_nl = for_equal_tmp_62 & (~ or_tmp_643);
  assign for_and_247_nl = for_equal_tmp_65 & (~ or_tmp_643);
  assign for_and_245_nl = for_equal_tmp_61 & (~ or_tmp_643);
  assign for_and_243_nl = for_equal_tmp_66 & (~ or_tmp_643);
  assign for_and_241_nl = for_equal_tmp_60 & (~ or_tmp_643);
  assign for_and_239_nl = for_equal_tmp_67 & (~ or_tmp_643);
  assign for_and_237_nl = for_equal_tmp_59 & (~ or_tmp_643);
  assign for_and_235_nl = for_equal_tmp_68 & (~ or_tmp_643);
  assign for_and_233_nl = for_equal_tmp_58 & (~ or_tmp_643);
  assign for_and_231_nl = for_equal_tmp_69 & (~ or_tmp_643);
  assign for_and_229_nl = for_equal_tmp_57 & (~ or_tmp_643);
  assign for_and_227_nl = for_equal_tmp_70 & (~ or_tmp_643);
  assign for_and_225_nl = for_equal_tmp_56 & (~ or_tmp_643);
  assign for_and_223_nl = for_equal_tmp_71 & (~ or_tmp_643);
  assign for_and_221_nl = for_equal_tmp_55 & (~ or_tmp_643);
  assign for_and_219_nl = for_equal_tmp_72 & (~ or_tmp_643);
  assign for_and_217_nl = for_equal_tmp_54 & (~ or_tmp_643);
  assign for_and_215_nl = for_equal_tmp_73 & (~ or_tmp_643);
  assign for_and_213_nl = for_equal_tmp_53 & (~ or_tmp_643);
  assign for_and_211_nl = for_equal_tmp_74 & (~ or_tmp_643);
  assign for_and_209_nl = for_equal_tmp_52 & (~ or_tmp_643);
  assign for_and_207_nl = for_equal_tmp_75 & (~ or_tmp_643);
  assign for_and_205_nl = for_equal_tmp_51 & (~ or_tmp_643);
  assign for_and_203_nl = for_equal_tmp_76 & (~ or_tmp_643);
  assign for_and_201_nl = for_equal_tmp_50 & (~ or_tmp_643);
  assign for_and_199_nl = for_equal_tmp_77 & (~ or_tmp_643);
  assign for_and_197_nl = for_equal_tmp_49 & (~ or_tmp_643);
  assign for_and_195_nl = for_equal_tmp_78 & (~ or_tmp_643);
  assign for_and_193_nl = for_equal_tmp_48 & (~ or_tmp_643);
  assign for_and_191_nl = for_equal_tmp_79 & (~ or_tmp_643);
  assign for_and_189_nl = for_equal_tmp_47 & (~ or_tmp_643);
  assign for_and_187_nl = for_equal_tmp_80 & (~ or_tmp_643);
  assign for_and_185_nl = for_equal_tmp_46 & (~ or_tmp_643);
  assign for_and_183_nl = for_equal_tmp_81 & (~ or_tmp_643);
  assign for_and_181_nl = for_equal_tmp_45 & (~ or_tmp_643);
  assign for_and_179_nl = for_equal_tmp_82 & (~ or_tmp_643);
  assign for_and_177_nl = for_equal_tmp_44 & (~ or_tmp_643);
  assign for_and_175_nl = for_equal_tmp_83 & (~ or_tmp_643);
  assign for_and_173_nl = for_equal_tmp_43 & (~ or_tmp_643);
  assign for_and_171_nl = for_equal_tmp_84 & (~ or_tmp_643);
  assign for_and_169_nl = for_equal_tmp_42 & (~ or_tmp_643);
  assign for_and_167_nl = for_equal_tmp_85 & (~ or_tmp_643);
  assign for_and_165_nl = for_equal_tmp_41 & (~ or_tmp_643);
  assign for_and_163_nl = for_equal_tmp_86 & (~ or_tmp_643);
  assign for_and_161_nl = for_equal_tmp_40 & (~ or_tmp_643);
  assign for_and_159_nl = for_equal_tmp_87 & (~ or_tmp_643);
  assign for_and_157_nl = for_equal_tmp_39 & (~ or_tmp_643);
  assign for_and_155_nl = for_equal_tmp_88 & (~ or_tmp_643);
  assign for_and_153_nl = for_equal_tmp_38 & (~ or_tmp_643);
  assign for_and_151_nl = for_equal_tmp_89 & (~ or_tmp_643);
  assign for_and_149_nl = for_equal_tmp_37 & (~ or_tmp_643);
  assign for_and_147_nl = for_equal_tmp_90 & (~ or_tmp_643);
  assign for_and_145_nl = for_equal_tmp_36 & (~ or_tmp_643);
  assign for_and_143_nl = for_equal_tmp_91 & (~ or_tmp_643);
  assign for_and_141_nl = for_equal_tmp_35 & (~ or_tmp_643);
  assign for_and_139_nl = for_equal_tmp_92 & (~ or_tmp_643);
  assign for_and_137_nl = for_equal_tmp_34 & (~ or_tmp_643);
  assign for_and_135_nl = for_equal_tmp_93 & (~ or_tmp_643);
  assign for_and_133_nl = for_equal_tmp_33 & (~ or_tmp_643);
  assign for_and_131_nl = for_equal_tmp_94 & (~ or_tmp_643);
  assign for_and_129_nl = or_dcpl_335 & (~ or_tmp_643);
  assign for_and_127_nl = for_equal_tmp_95 & (~ or_tmp_643);
  assign for_and_125_nl = for_equal_tmp_31 & (~ or_tmp_643);
  assign for_and_123_nl = for_equal_tmp_96 & (~ or_tmp_643);
  assign for_and_121_nl = for_equal_tmp_30 & (~ or_tmp_643);
  assign for_and_119_nl = for_equal_tmp_97 & (~ or_tmp_643);
  assign for_and_117_nl = for_equal_tmp_29 & (~ or_tmp_643);
  assign for_and_115_nl = for_equal_tmp_98 & (~ or_tmp_643);
  assign for_and_113_nl = for_equal_tmp_28 & (~ or_tmp_643);
  assign for_and_111_nl = for_equal_tmp_99 & (~ or_tmp_643);
  assign for_and_109_nl = for_equal_tmp_27 & (~ or_tmp_643);
  assign for_and_107_nl = for_equal_tmp_100 & (~ or_tmp_643);
  assign for_and_105_nl = for_equal_tmp_26 & (~ or_tmp_643);
  assign for_and_103_nl = for_equal_tmp_101 & (~ or_tmp_643);
  assign for_and_101_nl = for_equal_tmp_25 & (~ or_tmp_643);
  assign for_and_99_nl = for_equal_tmp_102 & (~ or_tmp_643);
  assign for_and_97_nl = for_equal_tmp_24 & (~ or_tmp_643);
  assign for_and_95_nl = for_equal_tmp_103 & (~ or_tmp_643);
  assign for_and_93_nl = for_equal_tmp_23 & (~ or_tmp_643);
  assign for_and_91_nl = for_equal_tmp_104 & (~ or_tmp_643);
  assign for_and_89_nl = for_equal_tmp_22 & (~ or_tmp_643);
  assign for_and_87_nl = for_equal_tmp_105 & (~ or_tmp_643);
  assign for_and_85_nl = for_equal_tmp_21 & (~ or_tmp_643);
  assign for_and_83_nl = for_equal_tmp_106 & (~ or_tmp_643);
  assign for_and_81_nl = for_equal_tmp_20 & (~ or_tmp_643);
  assign for_and_79_nl = for_equal_tmp_107 & (~ or_tmp_643);
  assign for_and_77_nl = for_equal_tmp_19 & (~ or_tmp_643);
  assign for_and_75_nl = for_equal_tmp_108 & (~ or_tmp_643);
  assign for_and_73_nl = for_equal_tmp_18 & (~ or_tmp_643);
  assign for_and_71_nl = for_equal_tmp_109 & (~ or_tmp_643);
  assign for_and_69_nl = for_equal_tmp_17 & (~ or_tmp_643);
  assign for_and_67_nl = for_equal_tmp_110 & (~ or_tmp_643);
  assign for_and_65_nl = or_dcpl_334 & (~ or_tmp_643);
  assign for_and_63_nl = for_equal_tmp_111 & (~ or_tmp_643);
  assign for_and_61_nl = for_equal_tmp_15 & (~ or_tmp_643);
  assign for_and_59_nl = for_equal_tmp_112 & (~ or_tmp_643);
  assign for_and_57_nl = for_equal_tmp_14 & (~ or_tmp_643);
  assign for_and_55_nl = for_equal_tmp_113 & (~ or_tmp_643);
  assign for_and_53_nl = for_equal_tmp_13 & (~ or_tmp_643);
  assign for_and_51_nl = for_equal_tmp_114 & (~ or_tmp_643);
  assign for_and_49_nl = for_equal_tmp_12 & (~ or_tmp_643);
  assign for_and_47_nl = for_equal_tmp_115 & (~ or_tmp_643);
  assign for_and_45_nl = for_equal_tmp_11 & (~ or_tmp_643);
  assign for_and_43_nl = for_equal_tmp_116 & (~ or_tmp_643);
  assign for_and_41_nl = for_equal_tmp_10 & (~ or_tmp_643);
  assign for_and_39_nl = for_equal_tmp_117 & (~ or_tmp_643);
  assign for_and_37_nl = for_equal_tmp_9 & (~ or_tmp_643);
  assign for_and_35_nl = for_equal_tmp_118 & (~ or_tmp_643);
  assign for_and_33_nl = or_dcpl_333 & (~ or_tmp_643);
  assign for_and_31_nl = for_equal_tmp_119 & (~ or_tmp_643);
  assign for_and_29_nl = for_equal_tmp_7 & (~ or_tmp_643);
  assign for_and_27_nl = for_equal_tmp_120 & (~ or_tmp_643);
  assign for_and_25_nl = for_equal_tmp_6 & (~ or_tmp_643);
  assign for_and_23_nl = for_equal_tmp_121 & (~ or_tmp_643);
  assign for_and_21_nl = for_equal_tmp_5 & (~ or_tmp_643);
  assign for_and_19_nl = for_equal_tmp_122 & (~ or_tmp_643);
  assign for_and_17_nl = or_dcpl_332 & (~ or_tmp_643);
  assign for_and_15_nl = for_equal_tmp_123 & (~ or_tmp_643);
  assign for_and_13_nl = for_equal_tmp_3 & (~ or_tmp_643);
  assign for_and_11_nl = for_equal_tmp_124 & (~ or_tmp_643);
  assign for_and_9_nl = or_dcpl_331 & (~ or_tmp_643);
  assign for_and_7_nl = for_equal_tmp_125 & (~ or_tmp_643);
  assign for_and_5_nl = or_dcpl_330 & (~ or_tmp_643);
  assign for_and_3_nl = for_equal_tmp_126 & (~ or_tmp_643);
  assign for_and_1_nl = for_equal_tmp_127 & (~ or_tmp_643);
  assign nl_i_7_0_sva_1  = conv_u2s_7_8(i_7_0_sva_6_0) + 8'b00000001;

  function automatic [31:0] MUX_v_32_128_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [31:0] input_3;
    input [31:0] input_4;
    input [31:0] input_5;
    input [31:0] input_6;
    input [31:0] input_7;
    input [31:0] input_8;
    input [31:0] input_9;
    input [31:0] input_10;
    input [31:0] input_11;
    input [31:0] input_12;
    input [31:0] input_13;
    input [31:0] input_14;
    input [31:0] input_15;
    input [31:0] input_16;
    input [31:0] input_17;
    input [31:0] input_18;
    input [31:0] input_19;
    input [31:0] input_20;
    input [31:0] input_21;
    input [31:0] input_22;
    input [31:0] input_23;
    input [31:0] input_24;
    input [31:0] input_25;
    input [31:0] input_26;
    input [31:0] input_27;
    input [31:0] input_28;
    input [31:0] input_29;
    input [31:0] input_30;
    input [31:0] input_31;
    input [31:0] input_32;
    input [31:0] input_33;
    input [31:0] input_34;
    input [31:0] input_35;
    input [31:0] input_36;
    input [31:0] input_37;
    input [31:0] input_38;
    input [31:0] input_39;
    input [31:0] input_40;
    input [31:0] input_41;
    input [31:0] input_42;
    input [31:0] input_43;
    input [31:0] input_44;
    input [31:0] input_45;
    input [31:0] input_46;
    input [31:0] input_47;
    input [31:0] input_48;
    input [31:0] input_49;
    input [31:0] input_50;
    input [31:0] input_51;
    input [31:0] input_52;
    input [31:0] input_53;
    input [31:0] input_54;
    input [31:0] input_55;
    input [31:0] input_56;
    input [31:0] input_57;
    input [31:0] input_58;
    input [31:0] input_59;
    input [31:0] input_60;
    input [31:0] input_61;
    input [31:0] input_62;
    input [31:0] input_63;
    input [31:0] input_64;
    input [31:0] input_65;
    input [31:0] input_66;
    input [31:0] input_67;
    input [31:0] input_68;
    input [31:0] input_69;
    input [31:0] input_70;
    input [31:0] input_71;
    input [31:0] input_72;
    input [31:0] input_73;
    input [31:0] input_74;
    input [31:0] input_75;
    input [31:0] input_76;
    input [31:0] input_77;
    input [31:0] input_78;
    input [31:0] input_79;
    input [31:0] input_80;
    input [31:0] input_81;
    input [31:0] input_82;
    input [31:0] input_83;
    input [31:0] input_84;
    input [31:0] input_85;
    input [31:0] input_86;
    input [31:0] input_87;
    input [31:0] input_88;
    input [31:0] input_89;
    input [31:0] input_90;
    input [31:0] input_91;
    input [31:0] input_92;
    input [31:0] input_93;
    input [31:0] input_94;
    input [31:0] input_95;
    input [31:0] input_96;
    input [31:0] input_97;
    input [31:0] input_98;
    input [31:0] input_99;
    input [31:0] input_100;
    input [31:0] input_101;
    input [31:0] input_102;
    input [31:0] input_103;
    input [31:0] input_104;
    input [31:0] input_105;
    input [31:0] input_106;
    input [31:0] input_107;
    input [31:0] input_108;
    input [31:0] input_109;
    input [31:0] input_110;
    input [31:0] input_111;
    input [31:0] input_112;
    input [31:0] input_113;
    input [31:0] input_114;
    input [31:0] input_115;
    input [31:0] input_116;
    input [31:0] input_117;
    input [31:0] input_118;
    input [31:0] input_119;
    input [31:0] input_120;
    input [31:0] input_121;
    input [31:0] input_122;
    input [31:0] input_123;
    input [31:0] input_124;
    input [31:0] input_125;
    input [31:0] input_126;
    input [31:0] input_127;
    input [6:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      7'b0000000 : begin
        result = input_0;
      end
      7'b0000001 : begin
        result = input_1;
      end
      7'b0000010 : begin
        result = input_2;
      end
      7'b0000011 : begin
        result = input_3;
      end
      7'b0000100 : begin
        result = input_4;
      end
      7'b0000101 : begin
        result = input_5;
      end
      7'b0000110 : begin
        result = input_6;
      end
      7'b0000111 : begin
        result = input_7;
      end
      7'b0001000 : begin
        result = input_8;
      end
      7'b0001001 : begin
        result = input_9;
      end
      7'b0001010 : begin
        result = input_10;
      end
      7'b0001011 : begin
        result = input_11;
      end
      7'b0001100 : begin
        result = input_12;
      end
      7'b0001101 : begin
        result = input_13;
      end
      7'b0001110 : begin
        result = input_14;
      end
      7'b0001111 : begin
        result = input_15;
      end
      7'b0010000 : begin
        result = input_16;
      end
      7'b0010001 : begin
        result = input_17;
      end
      7'b0010010 : begin
        result = input_18;
      end
      7'b0010011 : begin
        result = input_19;
      end
      7'b0010100 : begin
        result = input_20;
      end
      7'b0010101 : begin
        result = input_21;
      end
      7'b0010110 : begin
        result = input_22;
      end
      7'b0010111 : begin
        result = input_23;
      end
      7'b0011000 : begin
        result = input_24;
      end
      7'b0011001 : begin
        result = input_25;
      end
      7'b0011010 : begin
        result = input_26;
      end
      7'b0011011 : begin
        result = input_27;
      end
      7'b0011100 : begin
        result = input_28;
      end
      7'b0011101 : begin
        result = input_29;
      end
      7'b0011110 : begin
        result = input_30;
      end
      7'b0011111 : begin
        result = input_31;
      end
      7'b0100000 : begin
        result = input_32;
      end
      7'b0100001 : begin
        result = input_33;
      end
      7'b0100010 : begin
        result = input_34;
      end
      7'b0100011 : begin
        result = input_35;
      end
      7'b0100100 : begin
        result = input_36;
      end
      7'b0100101 : begin
        result = input_37;
      end
      7'b0100110 : begin
        result = input_38;
      end
      7'b0100111 : begin
        result = input_39;
      end
      7'b0101000 : begin
        result = input_40;
      end
      7'b0101001 : begin
        result = input_41;
      end
      7'b0101010 : begin
        result = input_42;
      end
      7'b0101011 : begin
        result = input_43;
      end
      7'b0101100 : begin
        result = input_44;
      end
      7'b0101101 : begin
        result = input_45;
      end
      7'b0101110 : begin
        result = input_46;
      end
      7'b0101111 : begin
        result = input_47;
      end
      7'b0110000 : begin
        result = input_48;
      end
      7'b0110001 : begin
        result = input_49;
      end
      7'b0110010 : begin
        result = input_50;
      end
      7'b0110011 : begin
        result = input_51;
      end
      7'b0110100 : begin
        result = input_52;
      end
      7'b0110101 : begin
        result = input_53;
      end
      7'b0110110 : begin
        result = input_54;
      end
      7'b0110111 : begin
        result = input_55;
      end
      7'b0111000 : begin
        result = input_56;
      end
      7'b0111001 : begin
        result = input_57;
      end
      7'b0111010 : begin
        result = input_58;
      end
      7'b0111011 : begin
        result = input_59;
      end
      7'b0111100 : begin
        result = input_60;
      end
      7'b0111101 : begin
        result = input_61;
      end
      7'b0111110 : begin
        result = input_62;
      end
      7'b0111111 : begin
        result = input_63;
      end
      7'b1000000 : begin
        result = input_64;
      end
      7'b1000001 : begin
        result = input_65;
      end
      7'b1000010 : begin
        result = input_66;
      end
      7'b1000011 : begin
        result = input_67;
      end
      7'b1000100 : begin
        result = input_68;
      end
      7'b1000101 : begin
        result = input_69;
      end
      7'b1000110 : begin
        result = input_70;
      end
      7'b1000111 : begin
        result = input_71;
      end
      7'b1001000 : begin
        result = input_72;
      end
      7'b1001001 : begin
        result = input_73;
      end
      7'b1001010 : begin
        result = input_74;
      end
      7'b1001011 : begin
        result = input_75;
      end
      7'b1001100 : begin
        result = input_76;
      end
      7'b1001101 : begin
        result = input_77;
      end
      7'b1001110 : begin
        result = input_78;
      end
      7'b1001111 : begin
        result = input_79;
      end
      7'b1010000 : begin
        result = input_80;
      end
      7'b1010001 : begin
        result = input_81;
      end
      7'b1010010 : begin
        result = input_82;
      end
      7'b1010011 : begin
        result = input_83;
      end
      7'b1010100 : begin
        result = input_84;
      end
      7'b1010101 : begin
        result = input_85;
      end
      7'b1010110 : begin
        result = input_86;
      end
      7'b1010111 : begin
        result = input_87;
      end
      7'b1011000 : begin
        result = input_88;
      end
      7'b1011001 : begin
        result = input_89;
      end
      7'b1011010 : begin
        result = input_90;
      end
      7'b1011011 : begin
        result = input_91;
      end
      7'b1011100 : begin
        result = input_92;
      end
      7'b1011101 : begin
        result = input_93;
      end
      7'b1011110 : begin
        result = input_94;
      end
      7'b1011111 : begin
        result = input_95;
      end
      7'b1100000 : begin
        result = input_96;
      end
      7'b1100001 : begin
        result = input_97;
      end
      7'b1100010 : begin
        result = input_98;
      end
      7'b1100011 : begin
        result = input_99;
      end
      7'b1100100 : begin
        result = input_100;
      end
      7'b1100101 : begin
        result = input_101;
      end
      7'b1100110 : begin
        result = input_102;
      end
      7'b1100111 : begin
        result = input_103;
      end
      7'b1101000 : begin
        result = input_104;
      end
      7'b1101001 : begin
        result = input_105;
      end
      7'b1101010 : begin
        result = input_106;
      end
      7'b1101011 : begin
        result = input_107;
      end
      7'b1101100 : begin
        result = input_108;
      end
      7'b1101101 : begin
        result = input_109;
      end
      7'b1101110 : begin
        result = input_110;
      end
      7'b1101111 : begin
        result = input_111;
      end
      7'b1110000 : begin
        result = input_112;
      end
      7'b1110001 : begin
        result = input_113;
      end
      7'b1110010 : begin
        result = input_114;
      end
      7'b1110011 : begin
        result = input_115;
      end
      7'b1110100 : begin
        result = input_116;
      end
      7'b1110101 : begin
        result = input_117;
      end
      7'b1110110 : begin
        result = input_118;
      end
      7'b1110111 : begin
        result = input_119;
      end
      7'b1111000 : begin
        result = input_120;
      end
      7'b1111001 : begin
        result = input_121;
      end
      7'b1111010 : begin
        result = input_122;
      end
      7'b1111011 : begin
        result = input_123;
      end
      7'b1111100 : begin
        result = input_124;
      end
      7'b1111101 : begin
        result = input_125;
      end
      7'b1111110 : begin
        result = input_126;
      end
      default : begin
        result = input_127;
      end
    endcase
    MUX_v_32_128_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [7:0] conv_u2s_7_8 ;
    input [6:0]  vector ;
  begin
    conv_u2s_7_8 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    fir
// ------------------------------------------------------------------


module fir (
  clk, rst, input_rsc_dat, input_rsc_triosy_lz, output_rsc_dat, output_rsc_triosy_lz
);
  input clk;
  input rst;
  input [4095:0] input_rsc_dat;
  output input_rsc_triosy_lz;
  output [4095:0] output_rsc_dat;
  output output_rsc_triosy_lz;



  // Interconnect Declarations for Component Instantiations 
  fir_core fir_core_inst (
      .clk(clk),
      .rst(rst),
      .input_rsc_dat(input_rsc_dat),
      .input_rsc_triosy_lz(input_rsc_triosy_lz),
      .output_rsc_dat(output_rsc_dat),
      .output_rsc_triosy_lz(output_rsc_triosy_lz)
    );
endmodule



